*Frequency Divide by 2 using E-TSPC Flip Flop
.include sky130nm.lib

xm1 1 out stage1 1 sky130_fd_pr__pfet_01v8 l=150n w=3050n 
xm2 stage1 clk 0 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm3 1 stage1 stage2 1 sky130_fd_pr__pfet_01v8 l=150n w=420n 
xm4 stage2 clk 0 0 sky130_fd_pr__nfet_01v8 l=150n w=840n

xm5 1 clk out 1 sky130_fd_pr__pfet_01v8 l=150n w=420n 
xm6 out stage2 0 0 sky130_fd_pr__nfet_01v8 l=150n w=840n

*output cap
c1 out 0 1f

*sources
v1 1 0 1.8
v2 clk 0 pulse(0 1.8 0 1ns 1ns 100ns 200ns)

*simulation
.control
tran 1ns 3us 400ns
plot v(clk)+2 v(out)
plot v(clk)+2 v(stage2)
plot v(clk)+2 v(stage1)
.endc
.end 
