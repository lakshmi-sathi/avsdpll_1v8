magic
tech sky130A
magscale 1 2
timestamp 1607692587
<< nwell >>
rect 178 1070 1534 1280
rect 274 958 1534 1070
rect 1010 920 1534 958
rect 1354 614 1534 616
rect 886 590 1534 614
rect 794 314 1534 590
rect 794 62 1028 314
<< pwell >>
rect 896 784 978 820
rect 896 694 978 730
<< nmos >>
rect 140 794 620 824
rect 140 682 500 712
rect 1108 712 1138 808
rect 1210 712 1240 808
rect 140 568 228 598
rect 398 172 428 256
rect 512 184 542 544
rect 624 184 654 664
rect 1158 142 1188 238
rect 1260 142 1290 238
<< pmos >>
rect 310 1060 440 1090
rect 574 1060 704 1090
rect 1108 1004 1138 1148
rect 1210 1004 1240 1148
rect 896 414 926 544
rect 1158 434 1188 578
rect 1260 434 1290 578
rect 896 150 926 280
<< ndiff >>
rect 140 874 620 890
rect 140 840 198 874
rect 232 840 266 874
rect 300 840 334 874
rect 368 840 402 874
rect 436 840 470 874
rect 504 840 538 874
rect 572 840 620 874
rect 140 824 620 840
rect 140 778 620 794
rect 1046 788 1108 808
rect 140 744 148 778
rect 182 744 216 778
rect 250 744 284 778
rect 318 744 352 778
rect 386 744 420 778
rect 454 744 522 778
rect 556 744 620 778
rect 140 730 620 744
rect 1046 754 1058 788
rect 1092 754 1108 788
rect 140 712 500 730
rect 140 616 500 682
rect 1046 712 1108 754
rect 1138 760 1210 808
rect 1138 726 1164 760
rect 1198 726 1210 760
rect 1138 712 1210 726
rect 1240 778 1298 808
rect 1240 744 1256 778
rect 1290 744 1298 778
rect 1240 712 1298 744
rect 560 634 624 664
rect 140 598 228 616
rect 560 600 574 634
rect 608 600 624 634
rect 140 552 228 568
rect 140 518 160 552
rect 194 518 228 552
rect 140 502 228 518
rect 560 566 624 600
rect 560 544 574 566
rect 446 256 512 544
rect 332 236 398 256
rect 332 202 348 236
rect 382 202 398 236
rect 332 172 398 202
rect 428 184 512 256
rect 542 532 574 544
rect 608 532 624 566
rect 542 498 624 532
rect 542 464 574 498
rect 608 464 624 498
rect 542 430 624 464
rect 542 396 574 430
rect 608 396 624 430
rect 542 362 624 396
rect 542 328 574 362
rect 608 328 624 362
rect 542 294 624 328
rect 542 260 574 294
rect 608 260 624 294
rect 542 226 624 260
rect 542 192 574 226
rect 608 192 624 226
rect 542 184 624 192
rect 654 602 720 664
rect 654 568 670 602
rect 704 568 720 602
rect 654 534 720 568
rect 654 500 670 534
rect 704 500 720 534
rect 654 430 720 500
rect 654 396 670 430
rect 704 396 720 430
rect 654 362 720 396
rect 654 328 670 362
rect 704 328 720 362
rect 654 294 720 328
rect 654 260 670 294
rect 704 260 720 294
rect 654 226 720 260
rect 654 192 670 226
rect 704 192 720 226
rect 654 184 720 192
rect 428 172 480 184
rect 1096 218 1158 238
rect 1096 184 1108 218
rect 1142 184 1158 218
rect 1096 142 1158 184
rect 1188 190 1260 238
rect 1188 156 1214 190
rect 1248 156 1260 190
rect 1188 142 1260 156
rect 1290 208 1348 238
rect 1290 174 1306 208
rect 1340 174 1348 208
rect 1290 142 1348 174
<< pdiff >>
rect 310 1140 440 1156
rect 310 1106 318 1140
rect 352 1106 386 1140
rect 420 1106 440 1140
rect 574 1140 704 1156
rect 310 1090 440 1106
rect 310 1044 440 1060
rect 310 1010 326 1044
rect 360 1010 398 1044
rect 432 1010 440 1044
rect 574 1106 582 1140
rect 616 1106 650 1140
rect 684 1106 704 1140
rect 574 1090 704 1106
rect 1046 1140 1108 1148
rect 1046 1106 1058 1140
rect 1092 1106 1108 1140
rect 1046 1072 1108 1106
rect 574 1044 704 1060
rect 310 994 440 1010
rect 574 1010 592 1044
rect 626 1010 660 1044
rect 694 1010 704 1044
rect 574 994 704 1010
rect 1046 1038 1058 1072
rect 1092 1038 1108 1072
rect 1046 1004 1108 1038
rect 1138 1140 1210 1148
rect 1138 1106 1164 1140
rect 1198 1106 1210 1140
rect 1138 1072 1210 1106
rect 1138 1038 1164 1072
rect 1198 1038 1210 1072
rect 1138 1004 1210 1038
rect 1240 1140 1300 1148
rect 1240 1106 1254 1140
rect 1288 1106 1300 1140
rect 1240 1072 1300 1106
rect 1240 1038 1254 1072
rect 1288 1038 1300 1072
rect 1240 1004 1300 1038
rect 1096 570 1158 578
rect 830 534 896 544
rect 830 500 846 534
rect 880 500 896 534
rect 830 466 896 500
rect 830 432 846 466
rect 880 432 896 466
rect 830 414 896 432
rect 926 524 992 544
rect 926 490 942 524
rect 976 490 992 524
rect 926 456 992 490
rect 926 422 942 456
rect 976 422 992 456
rect 1096 536 1108 570
rect 1142 536 1158 570
rect 1096 502 1158 536
rect 1096 468 1108 502
rect 1142 468 1158 502
rect 1096 434 1158 468
rect 1188 570 1260 578
rect 1188 536 1214 570
rect 1248 536 1260 570
rect 1188 502 1260 536
rect 1188 468 1214 502
rect 1248 468 1260 502
rect 1188 434 1260 468
rect 1290 570 1350 578
rect 1290 536 1304 570
rect 1338 536 1350 570
rect 1290 502 1350 536
rect 1290 468 1304 502
rect 1338 468 1350 502
rect 1290 434 1350 468
rect 926 414 992 422
rect 830 272 896 280
rect 830 238 846 272
rect 880 238 896 272
rect 830 200 896 238
rect 830 166 846 200
rect 880 166 896 200
rect 830 150 896 166
rect 926 260 992 280
rect 926 226 942 260
rect 976 226 992 260
rect 926 192 992 226
rect 926 158 942 192
rect 976 158 992 192
rect 926 150 992 158
<< ndiffc >>
rect 198 840 232 874
rect 266 840 300 874
rect 334 840 368 874
rect 402 840 436 874
rect 470 840 504 874
rect 538 840 572 874
rect 148 744 182 778
rect 216 744 250 778
rect 284 744 318 778
rect 352 744 386 778
rect 420 744 454 778
rect 522 744 556 778
rect 1058 754 1092 788
rect 1164 726 1198 760
rect 1256 744 1290 778
rect 574 600 608 634
rect 160 518 194 552
rect 348 202 382 236
rect 574 532 608 566
rect 574 464 608 498
rect 574 396 608 430
rect 574 328 608 362
rect 574 260 608 294
rect 574 192 608 226
rect 670 568 704 602
rect 670 500 704 534
rect 670 396 704 430
rect 670 328 704 362
rect 670 260 704 294
rect 670 192 704 226
rect 1108 184 1142 218
rect 1214 156 1248 190
rect 1306 174 1340 208
<< pdiffc >>
rect 318 1106 352 1140
rect 386 1106 420 1140
rect 326 1010 360 1044
rect 398 1010 432 1044
rect 582 1106 616 1140
rect 650 1106 684 1140
rect 1058 1106 1092 1140
rect 592 1010 626 1044
rect 660 1010 694 1044
rect 1058 1038 1092 1072
rect 1164 1106 1198 1140
rect 1164 1038 1198 1072
rect 1254 1106 1288 1140
rect 1254 1038 1288 1072
rect 846 500 880 534
rect 846 432 880 466
rect 942 490 976 524
rect 942 422 976 456
rect 1108 536 1142 570
rect 1108 468 1142 502
rect 1214 536 1248 570
rect 1214 468 1248 502
rect 1304 536 1338 570
rect 1304 468 1338 502
rect 846 238 880 272
rect 846 166 880 200
rect 942 226 976 260
rect 942 158 976 192
<< psubdiff >>
rect 896 786 920 820
rect 954 786 978 820
rect 896 784 978 786
rect 896 696 920 730
rect 954 696 978 730
rect 896 694 978 696
<< nsubdiff >>
rect 228 1210 256 1244
rect 290 1210 314 1244
rect 392 1210 420 1244
rect 454 1210 478 1244
rect 558 1210 584 1244
rect 618 1210 642 1244
rect 718 1210 748 1244
rect 782 1210 806 1244
rect 886 1210 912 1244
rect 946 1210 970 1244
rect 1406 536 1432 570
rect 1466 536 1492 570
rect 1406 534 1492 536
rect 1406 478 1492 480
rect 1406 444 1432 478
rect 1466 444 1492 478
rect 1406 442 1492 444
rect 1406 386 1492 388
rect 1406 352 1432 386
rect 1466 352 1492 386
rect 1406 350 1492 352
<< psubdiffcont >>
rect 920 786 954 820
rect 920 696 954 730
<< nsubdiffcont >>
rect 256 1210 290 1244
rect 420 1210 454 1244
rect 584 1210 618 1244
rect 748 1210 782 1244
rect 912 1210 946 1244
rect 1432 536 1466 570
rect 1432 444 1466 478
rect 1432 352 1466 386
<< poly >>
rect 1108 1148 1138 1174
rect 1210 1148 1240 1174
rect 480 1092 534 1108
rect 480 1090 490 1092
rect 284 1060 310 1090
rect 440 1060 490 1090
rect 480 1058 490 1060
rect 524 1090 534 1092
rect 524 1060 574 1090
rect 704 1060 730 1090
rect 524 1058 534 1060
rect 480 1042 534 1058
rect 490 948 524 1042
rect 490 918 680 948
rect 1108 924 1138 1004
rect 1210 936 1240 1004
rect 646 824 680 918
rect 1082 914 1138 924
rect 1204 922 1240 936
rect 1076 880 1092 914
rect 1126 880 1140 914
rect 1182 904 1240 922
rect 1082 870 1138 880
rect 92 794 140 824
rect 620 794 680 824
rect 92 712 122 794
rect 1108 808 1138 870
rect 1182 870 1192 904
rect 1226 870 1240 904
rect 1182 854 1240 870
rect 1204 842 1240 854
rect 1210 808 1240 842
rect 16 686 140 712
rect 16 652 26 686
rect 60 682 140 686
rect 500 682 526 712
rect 60 652 70 682
rect 16 636 70 652
rect 624 680 788 712
rect 1108 686 1138 712
rect 1210 686 1240 712
rect 624 664 654 680
rect 114 568 140 598
rect 228 568 542 598
rect 248 562 542 568
rect 248 456 278 562
rect 512 544 542 562
rect 180 446 278 456
rect 180 412 196 446
rect 230 412 278 446
rect 180 402 278 412
rect 352 336 428 346
rect 352 302 368 336
rect 402 302 428 336
rect 352 292 428 302
rect 398 256 428 292
rect 748 364 788 680
rect 1158 578 1188 604
rect 1260 578 1290 604
rect 896 544 926 570
rect 896 374 926 414
rect 878 364 944 374
rect 748 330 894 364
rect 928 330 944 364
rect 1158 354 1188 434
rect 1260 366 1290 434
rect 1132 344 1188 354
rect 1254 352 1290 366
rect 878 320 944 330
rect 896 280 926 320
rect 1126 310 1142 344
rect 1176 310 1190 344
rect 1232 334 1290 352
rect 1132 300 1188 310
rect 398 146 428 172
rect 512 166 542 184
rect 624 166 654 184
rect 512 136 654 166
rect 1158 238 1188 300
rect 1232 300 1242 334
rect 1276 300 1290 334
rect 1232 284 1290 300
rect 1254 272 1290 284
rect 1260 238 1290 272
rect 896 124 926 150
rect 1158 116 1188 142
rect 1260 116 1290 142
<< polycont >>
rect 490 1058 524 1092
rect 1092 880 1126 914
rect 1192 870 1226 904
rect 26 652 60 686
rect 196 412 230 446
rect 368 302 402 336
rect 894 330 928 364
rect 1142 310 1176 344
rect 1242 300 1276 334
<< locali >>
rect 0 1210 160 1244
rect 194 1210 256 1244
rect 290 1210 296 1244
rect 330 1210 420 1244
rect 466 1210 568 1244
rect 618 1210 704 1244
rect 738 1210 748 1244
rect 782 1210 840 1244
rect 874 1210 912 1244
rect 946 1210 976 1244
rect 1010 1210 1112 1244
rect 1146 1210 1248 1244
rect 1282 1210 1534 1244
rect 330 1144 414 1210
rect 302 1140 444 1144
rect 302 1106 318 1140
rect 352 1106 386 1140
rect 420 1106 444 1140
rect 302 1102 444 1106
rect 484 1140 704 1142
rect 484 1106 582 1140
rect 616 1106 650 1140
rect 684 1106 704 1140
rect 484 1104 704 1106
rect 1052 1140 1096 1156
rect 1052 1106 1058 1140
rect 1092 1106 1096 1140
rect 484 1092 530 1104
rect 484 1058 490 1092
rect 524 1058 530 1092
rect 310 1044 448 1048
rect 310 1010 326 1044
rect 360 1010 398 1044
rect 432 1010 448 1044
rect 484 1042 530 1058
rect 1052 1072 1096 1106
rect 568 1044 710 1046
rect 310 976 448 1010
rect 74 926 448 976
rect 568 1010 592 1044
rect 626 1010 660 1044
rect 694 1010 710 1044
rect 568 1008 710 1010
rect 1052 1038 1058 1072
rect 1092 1038 1096 1072
rect 74 790 128 926
rect 568 914 656 1008
rect 1052 982 1096 1038
rect 1154 1140 1200 1210
rect 1154 1106 1164 1140
rect 1198 1106 1200 1140
rect 1154 1072 1200 1106
rect 1154 1038 1164 1072
rect 1198 1038 1200 1072
rect 1154 1016 1200 1038
rect 1254 1140 1312 1156
rect 1288 1106 1312 1140
rect 1254 1072 1312 1106
rect 1288 1038 1312 1072
rect 1254 1004 1312 1038
rect 1052 948 1220 982
rect 1180 922 1220 948
rect 568 890 1092 914
rect 174 880 1092 890
rect 1126 880 1142 914
rect 1180 904 1226 922
rect 174 874 658 880
rect 174 840 198 874
rect 232 840 266 874
rect 300 840 334 874
rect 368 840 402 874
rect 436 840 470 874
rect 504 840 538 874
rect 572 840 658 874
rect 1180 870 1192 904
rect 1180 854 1226 870
rect 1278 896 1312 1004
rect 1278 862 1630 896
rect 1180 846 1218 854
rect 174 838 658 840
rect 74 778 620 790
rect 74 744 148 778
rect 182 744 216 778
rect 250 744 284 778
rect 318 744 352 778
rect 386 744 420 778
rect 454 744 522 778
rect 556 744 620 778
rect 74 742 620 744
rect 868 786 920 820
rect 954 786 1002 820
rect 868 730 1002 786
rect 1050 812 1218 846
rect 1050 788 1094 812
rect 1278 808 1312 862
rect 1050 754 1058 788
rect 1092 754 1094 788
rect 1252 778 1312 808
rect 1050 736 1094 754
rect 1156 760 1200 776
rect 8 686 62 702
rect 8 652 26 686
rect 60 652 62 686
rect 868 696 920 730
rect 954 696 1002 730
rect 8 348 62 652
rect 572 634 610 664
rect 572 600 574 634
rect 608 600 610 634
rect 572 566 610 600
rect 156 552 198 556
rect 140 518 160 552
rect 194 518 212 552
rect 572 532 574 566
rect 608 532 610 566
rect 156 502 198 518
rect 572 498 610 532
rect 572 464 574 498
rect 608 464 610 498
rect 180 412 196 446
rect 230 412 246 446
rect 572 430 610 464
rect 572 396 574 430
rect 608 396 610 430
rect 572 362 610 396
rect -316 336 420 348
rect -316 302 368 336
rect 402 302 420 336
rect -316 290 420 302
rect 572 328 574 362
rect 608 328 610 362
rect 572 294 610 328
rect 346 236 382 256
rect 346 202 348 236
rect 346 184 382 202
rect 572 248 574 294
rect 608 248 610 294
rect 572 226 610 248
rect 572 192 574 226
rect 608 192 610 226
rect 572 172 610 192
rect 668 602 706 664
rect 868 658 1002 696
rect 1156 726 1164 760
rect 1198 726 1200 760
rect 1156 672 1200 726
rect 1252 744 1256 778
rect 1290 744 1312 778
rect 1252 712 1312 744
rect 1112 658 1246 672
rect 868 624 988 658
rect 1022 624 1124 658
rect 1158 624 1260 658
rect 1294 624 1534 658
rect 668 568 670 602
rect 704 568 706 602
rect 668 534 706 568
rect 1102 570 1146 586
rect 668 500 670 534
rect 704 502 706 534
rect 844 534 882 550
rect 844 524 846 534
rect 790 502 846 524
rect 704 500 846 502
rect 880 500 882 534
rect 668 480 882 500
rect 668 446 686 480
rect 720 466 882 480
rect 720 452 846 466
rect 720 446 728 452
rect 668 440 728 446
rect 668 430 720 440
rect 790 436 846 452
rect 668 396 670 430
rect 704 396 720 430
rect 844 432 846 436
rect 880 432 882 466
rect 844 414 882 432
rect 940 524 978 544
rect 940 490 942 524
rect 976 490 978 524
rect 940 456 978 490
rect 940 422 942 456
rect 976 422 978 456
rect 668 362 720 396
rect 940 370 978 422
rect 1102 536 1108 570
rect 1142 536 1146 570
rect 1102 502 1146 536
rect 1102 468 1108 502
rect 1142 468 1146 502
rect 1102 412 1146 468
rect 1204 570 1250 586
rect 1204 536 1214 570
rect 1248 536 1250 570
rect 1204 508 1250 536
rect 1304 570 1362 586
rect 1338 536 1362 570
rect 1204 502 1266 508
rect 1204 468 1214 502
rect 1248 496 1266 502
rect 1204 462 1232 468
rect 1204 450 1266 462
rect 1304 502 1362 536
rect 1406 536 1432 570
rect 1466 536 1492 570
rect 1406 534 1492 536
rect 1338 468 1362 502
rect 1420 480 1480 534
rect 1204 446 1250 450
rect 1102 378 1270 412
rect 1304 386 1362 468
rect 1406 478 1492 480
rect 1406 442 1432 478
rect 1420 441 1432 442
rect 1466 442 1492 478
rect 1466 441 1480 442
rect 1420 388 1480 441
rect 668 328 670 362
rect 704 328 720 362
rect 668 294 720 328
rect 878 364 978 370
rect 878 330 894 364
rect 928 330 978 364
rect 1232 352 1270 378
rect 878 324 978 330
rect 1028 310 1040 344
rect 1074 310 1142 344
rect 1176 310 1192 344
rect 1232 334 1276 352
rect 1232 300 1242 334
rect 1232 294 1276 300
rect 668 260 670 294
rect 704 260 720 294
rect 668 226 720 260
rect 668 192 670 226
rect 704 218 720 226
rect 792 272 884 288
rect 1230 284 1276 294
rect 792 238 846 272
rect 880 238 884 272
rect 792 234 884 238
rect 704 192 706 218
rect 668 172 706 192
rect 792 200 818 234
rect 852 200 884 234
rect 792 166 846 200
rect 880 166 884 200
rect 792 150 884 166
rect 938 260 980 284
rect 1230 276 1266 284
rect 938 226 942 260
rect 976 226 980 260
rect 938 192 980 226
rect 938 158 942 192
rect 976 158 980 192
rect 1100 242 1266 276
rect 1328 280 1362 386
rect 1406 386 1492 388
rect 1406 352 1432 386
rect 1466 352 1492 386
rect 1406 350 1492 352
rect 1328 246 1658 280
rect 1100 218 1144 242
rect 1328 238 1362 246
rect 1100 184 1108 218
rect 1142 184 1144 218
rect 1302 208 1362 238
rect 1100 166 1144 184
rect 1206 190 1250 206
rect 938 62 980 158
rect 1206 156 1214 190
rect 1248 156 1250 190
rect 1206 140 1250 156
rect 1302 174 1306 208
rect 1340 174 1362 208
rect 1302 142 1362 174
rect 0 28 160 62
rect 194 28 296 62
rect 330 28 432 62
rect 466 28 568 62
rect 602 28 704 62
rect 738 28 840 62
rect 874 28 976 62
rect 1010 28 1112 62
rect 1146 28 1248 62
rect 1282 28 1534 62
<< viali >>
rect 160 1210 194 1244
rect 296 1210 330 1244
rect 432 1210 454 1244
rect 454 1210 466 1244
rect 568 1210 584 1244
rect 584 1210 602 1244
rect 704 1210 738 1244
rect 840 1210 874 1244
rect 976 1210 1010 1244
rect 1112 1210 1146 1244
rect 1248 1210 1282 1244
rect 160 518 194 552
rect 196 412 230 446
rect 348 202 382 236
rect 574 260 608 282
rect 574 248 608 260
rect 988 624 1022 658
rect 1124 624 1158 658
rect 1260 624 1294 658
rect 686 446 720 480
rect 1232 468 1248 496
rect 1248 468 1266 496
rect 1232 462 1266 468
rect 1432 444 1466 475
rect 1432 441 1466 444
rect 1040 310 1074 344
rect 818 200 852 234
rect 1214 156 1248 190
rect 160 28 194 62
rect 296 28 330 62
rect 432 28 466 62
rect 568 28 602 62
rect 704 28 738 62
rect 840 28 874 62
rect 976 28 1010 62
rect 1112 28 1146 62
rect 1248 28 1282 62
<< metal1 >>
rect 0 1244 1534 1280
rect 0 1210 160 1244
rect 194 1210 296 1244
rect 330 1210 432 1244
rect 466 1210 568 1244
rect 602 1210 704 1244
rect 738 1210 840 1244
rect 874 1210 976 1244
rect 1010 1210 1112 1244
rect 1146 1210 1248 1244
rect 1282 1210 1534 1244
rect 0 1184 1534 1210
rect 0 658 1534 688
rect 0 624 988 658
rect 1022 624 1124 658
rect 1158 624 1260 658
rect 1294 624 1534 658
rect 0 592 1534 624
rect 148 552 208 592
rect 148 518 160 552
rect 194 518 208 552
rect 148 506 208 518
rect -340 446 242 458
rect -340 412 196 446
rect 230 412 242 446
rect -340 404 242 412
rect 142 402 242 404
rect 456 248 504 592
rect 668 489 738 498
rect 668 437 677 489
rect 729 437 738 489
rect 668 428 738 437
rect 1026 352 1090 358
rect 1026 300 1032 352
rect 1084 300 1090 352
rect 1026 294 1090 300
rect 336 236 504 248
rect 562 282 758 294
rect 562 248 574 282
rect 608 248 758 282
rect 562 246 758 248
rect 562 236 864 246
rect 336 202 348 236
rect 382 202 504 236
rect 336 190 504 202
rect 712 234 864 236
rect 712 200 818 234
rect 852 200 864 234
rect 712 188 864 200
rect 1120 202 1174 592
rect 1220 496 1482 508
rect 1220 462 1232 496
rect 1266 475 1482 496
rect 1266 462 1432 475
rect 1220 450 1432 462
rect 1312 441 1432 450
rect 1466 441 1482 475
rect 1312 414 1482 441
rect 1120 190 1254 202
rect 1120 156 1214 190
rect 1248 156 1254 190
rect 1120 144 1254 156
rect 1312 96 1372 414
rect 0 62 1534 96
rect 0 28 160 62
rect 194 28 296 62
rect 330 28 432 62
rect 466 28 568 62
rect 602 28 704 62
rect 738 28 840 62
rect 874 28 976 62
rect 1010 28 1112 62
rect 1146 28 1248 62
rect 1282 28 1534 62
rect 0 0 1534 28
<< via1 >>
rect 677 480 729 489
rect 677 446 686 480
rect 686 446 720 480
rect 720 446 729 480
rect 677 437 729 446
rect 1032 344 1084 352
rect 1032 310 1040 344
rect 1040 310 1074 344
rect 1074 310 1084 344
rect 1032 300 1084 310
<< metal2 >>
rect 668 492 738 498
rect 668 489 1080 492
rect 668 437 677 489
rect 729 438 1080 489
rect 729 437 738 438
rect 668 428 738 437
rect 1028 358 1080 438
rect 1026 352 1090 358
rect 1026 300 1032 352
rect 1084 300 1090 352
rect 1026 294 1090 300
<< labels >>
rlabel locali s 174 292 228 346 4 Clk_Ref
port 1 nsew
rlabel locali s 1278 866 1312 900 4 Up
port 2 nsew
rlabel locali s 1328 298 1362 332 4 Down
port 3 nsew
rlabel metal1 s 142 430 142 430 4 Clk2
port 4 nsew
rlabel metal1 s 0 640 0 640 4 GND
port 5 nsew
rlabel metal1 s 0 1232 0 1232 4 VDD
port 6 nsew
rlabel metal1 s 0 48 0 48 4 VDD
port 6 nsew
<< end >>
