magic
tech sky130A
timestamp 1605105670
<< nwell >>
rect -140 283 437 284
rect -140 171 539 283
rect -132 64 539 171
<< nmos >>
rect -83 -10 -68 26
rect 29 -10 44 26
rect 136 -55 151 29
rect 245 -10 260 26
rect 352 -55 367 29
rect 477 -10 492 26
<< pmos >>
rect -83 88 -68 160
rect 29 88 44 160
rect 136 82 151 124
rect 245 88 260 160
rect 352 82 367 124
rect 477 88 492 160
<< ndiff >>
rect -112 17 -83 26
rect -112 0 -106 17
rect -89 0 -83 17
rect -112 -10 -83 0
rect -68 17 -39 26
rect -68 0 -62 17
rect -45 0 -39 17
rect -68 -10 -39 0
rect 0 17 29 26
rect 0 0 6 17
rect 23 0 29 17
rect 0 -10 29 0
rect 44 17 73 26
rect 44 0 50 17
rect 67 0 73 17
rect 44 -10 73 0
rect 107 20 136 29
rect 107 3 113 20
rect 130 3 136 20
rect 107 -14 136 3
rect 107 -31 113 -14
rect 130 -31 136 -14
rect 107 -55 136 -31
rect 151 20 180 29
rect 151 3 157 20
rect 174 3 180 20
rect 151 -14 180 3
rect 216 17 245 26
rect 216 0 222 17
rect 239 0 245 17
rect 216 -10 245 0
rect 260 17 289 26
rect 260 0 266 17
rect 283 0 289 17
rect 260 -10 289 0
rect 323 20 352 29
rect 323 3 329 20
rect 346 3 352 20
rect 151 -31 157 -14
rect 174 -31 180 -14
rect 323 -14 352 3
rect 323 -31 329 -14
rect 346 -31 352 -14
rect 151 -55 180 -31
rect 323 -55 352 -31
rect 367 20 396 29
rect 367 3 373 20
rect 390 3 396 20
rect 367 -14 396 3
rect 448 17 477 26
rect 448 0 454 17
rect 471 0 477 17
rect 448 -10 477 0
rect 492 17 521 26
rect 492 0 498 17
rect 515 0 521 17
rect 492 -10 521 0
rect 367 -31 373 -14
rect 390 -31 396 -14
rect 367 -55 396 -31
<< pdiff >>
rect -112 156 -83 160
rect -112 139 -106 156
rect -89 139 -83 156
rect -112 122 -83 139
rect -112 105 -106 122
rect -89 105 -83 122
rect -112 88 -83 105
rect -68 143 -39 160
rect -68 126 -62 143
rect -45 126 -39 143
rect -68 109 -39 126
rect -68 92 -62 109
rect -45 92 -39 109
rect -68 88 -39 92
rect 0 156 29 160
rect 0 139 6 156
rect 23 139 29 156
rect 0 122 29 139
rect 0 105 6 122
rect 23 105 29 122
rect 0 88 29 105
rect 44 143 73 160
rect 44 126 50 143
rect 67 126 73 143
rect 44 109 73 126
rect 216 156 245 160
rect 216 139 222 156
rect 239 139 245 156
rect 44 92 50 109
rect 67 92 73 109
rect 44 88 73 92
rect 107 111 136 124
rect 107 94 113 111
rect 130 94 136 111
rect 107 82 136 94
rect 151 110 180 124
rect 151 93 157 110
rect 174 93 180 110
rect 151 82 180 93
rect 216 122 245 139
rect 216 105 222 122
rect 239 105 245 122
rect 216 88 245 105
rect 260 143 289 160
rect 448 156 477 160
rect 260 126 266 143
rect 283 126 289 143
rect 260 109 289 126
rect 448 139 454 156
rect 471 139 477 156
rect 260 92 266 109
rect 283 92 289 109
rect 260 88 289 92
rect 323 111 352 124
rect 323 94 329 111
rect 346 94 352 111
rect 323 82 352 94
rect 367 110 396 124
rect 367 93 373 110
rect 390 93 396 110
rect 367 82 396 93
rect 448 122 477 139
rect 448 105 454 122
rect 471 105 477 122
rect 448 88 477 105
rect 492 143 521 160
rect 492 126 498 143
rect 515 126 521 143
rect 492 109 521 126
rect 492 92 498 109
rect 515 92 521 109
rect 492 88 521 92
<< ndiffc >>
rect -106 0 -89 17
rect -62 0 -45 17
rect 6 0 23 17
rect 50 0 67 17
rect 113 3 130 20
rect 113 -31 130 -14
rect 157 3 174 20
rect 222 0 239 17
rect 266 0 283 17
rect 329 3 346 20
rect 157 -31 174 -14
rect 329 -31 346 -14
rect 373 3 390 20
rect 454 0 471 17
rect 498 0 515 17
rect 373 -31 390 -14
<< pdiffc >>
rect -106 139 -89 156
rect -106 105 -89 122
rect -62 126 -45 143
rect -62 92 -45 109
rect 6 139 23 156
rect 6 105 23 122
rect 50 126 67 143
rect 222 139 239 156
rect 50 92 67 109
rect 113 94 130 111
rect 157 93 174 110
rect 222 105 239 122
rect 266 126 283 143
rect 454 139 471 156
rect 266 92 283 109
rect 329 94 346 111
rect 373 93 390 110
rect 454 105 471 122
rect 498 126 515 143
rect 498 92 515 109
<< psubdiff >>
rect -123 -108 -110 -91
rect -93 -108 -81 -91
rect -39 -108 -26 -91
rect -9 -108 3 -91
rect 45 -108 58 -91
rect 75 -108 87 -91
rect 129 -108 142 -91
rect 159 -108 171 -91
rect 213 -108 226 -91
rect 243 -108 255 -91
rect 297 -108 310 -91
rect 327 -108 339 -91
rect 381 -108 394 -91
rect 411 -108 423 -91
rect 465 -108 478 -91
rect 495 -108 507 -91
<< nsubdiff >>
rect -114 246 -102 265
rect -83 246 -71 265
rect -28 246 -16 265
rect 3 246 15 265
rect 58 246 70 265
rect 89 246 101 265
rect 144 246 156 265
rect 175 246 187 265
rect 230 246 242 265
rect 261 246 273 265
rect 316 246 328 265
rect 347 246 359 265
rect 402 246 414 265
rect 433 246 445 265
<< psubdiffcont >>
rect -110 -108 -93 -91
rect -26 -108 -9 -91
rect 58 -108 75 -91
rect 142 -108 159 -91
rect 226 -108 243 -91
rect 310 -108 327 -91
rect 394 -108 411 -91
rect 478 -108 495 -91
<< nsubdiffcont >>
rect -102 246 -83 265
rect -16 246 3 265
rect 70 246 89 265
rect 156 246 175 265
rect 242 246 261 265
rect 328 246 347 265
rect 414 246 433 265
<< poly >>
rect 131 198 158 206
rect 131 181 136 198
rect 153 181 158 198
rect 131 173 158 181
rect -83 160 -68 173
rect 29 160 44 173
rect 136 124 151 173
rect 245 160 260 173
rect 347 169 380 174
rect -83 68 -68 88
rect 29 68 44 88
rect 347 152 355 169
rect 372 152 380 169
rect 477 160 492 173
rect 347 147 380 152
rect 352 124 367 147
rect 136 68 151 82
rect 245 68 260 88
rect 352 68 367 82
rect 477 68 492 88
rect -112 66 -68 68
rect 0 66 44 68
rect 216 66 260 68
rect 448 66 492 68
rect -115 63 -68 66
rect -115 46 -106 63
rect -89 46 -68 63
rect -115 42 -68 46
rect -3 63 44 66
rect -3 46 6 63
rect 23 46 44 63
rect -3 42 44 46
rect 213 63 260 66
rect 213 46 222 63
rect 239 46 260 63
rect 213 42 260 46
rect 445 63 492 66
rect 445 46 454 63
rect 471 46 492 63
rect 445 42 492 46
rect -112 41 -68 42
rect 0 41 44 42
rect -83 26 -68 41
rect 29 26 44 41
rect 136 29 151 42
rect 216 41 260 42
rect -83 -23 -68 -10
rect 29 -23 44 -10
rect 65 -29 92 -21
rect 65 -46 70 -29
rect 87 -46 92 -29
rect 65 -64 92 -46
rect 245 26 260 41
rect 352 29 367 42
rect 448 41 492 42
rect 245 -23 260 -10
rect 282 -40 309 -31
rect 136 -64 151 -55
rect 65 -81 151 -64
rect 282 -57 287 -40
rect 304 -57 309 -40
rect 477 26 492 41
rect 477 -23 492 -10
rect 282 -65 309 -57
rect 352 -65 367 -55
rect 282 -80 367 -65
<< polycont >>
rect 136 181 153 198
rect 355 152 372 169
rect -106 46 -89 63
rect 6 46 23 63
rect 222 46 239 63
rect 454 46 471 63
rect 70 -46 87 -29
rect 287 -57 304 -40
<< locali >>
rect -146 265 553 284
rect -146 246 -102 265
rect -83 246 -16 265
rect 3 246 70 265
rect 89 246 156 265
rect 175 246 242 265
rect 261 246 328 265
rect 347 246 414 265
rect 433 246 553 265
rect -146 236 553 246
rect -106 156 -89 236
rect -106 122 -89 139
rect -106 88 -89 105
rect -62 143 -45 160
rect -62 109 -45 126
rect -62 71 -45 92
rect 6 156 23 236
rect 136 214 153 218
rect 136 171 153 181
rect 6 122 23 139
rect 6 88 23 105
rect 50 143 67 160
rect 50 109 67 126
rect 222 156 239 236
rect 393 235 471 236
rect 50 71 67 92
rect 113 111 130 124
rect 113 71 130 94
rect -62 64 -32 71
rect -144 46 -106 63
rect -89 46 -81 63
rect -62 47 -56 64
rect -39 47 -32 64
rect -62 41 -32 47
rect -3 46 6 63
rect 23 46 31 63
rect 50 41 130 71
rect -106 17 -89 26
rect -106 -78 -89 0
rect -62 17 -45 41
rect -62 -10 -45 0
rect 6 17 23 26
rect 6 -49 23 0
rect 50 17 67 41
rect 50 -10 67 0
rect 113 20 130 41
rect 113 -14 130 3
rect 62 -46 70 -29
rect 87 -46 95 -29
rect 113 -39 130 -31
rect 157 110 174 124
rect 157 68 174 93
rect 222 122 239 139
rect 222 88 239 105
rect 266 143 283 160
rect 346 152 355 169
rect 372 152 380 169
rect 454 156 471 235
rect 266 109 283 126
rect 266 71 283 92
rect 329 111 346 124
rect 329 71 346 94
rect 157 63 243 68
rect 157 46 222 63
rect 239 46 247 63
rect 157 43 243 46
rect 157 20 174 43
rect 266 41 346 71
rect 157 -14 174 3
rect 157 -39 174 -31
rect 222 17 239 26
rect 5 -78 23 -49
rect 222 -51 239 0
rect 266 17 283 41
rect 266 -10 283 0
rect 329 20 346 41
rect 329 -14 346 3
rect 222 -78 240 -51
rect 271 -57 281 -36
rect 302 -37 307 -36
rect 302 -40 312 -37
rect 329 -39 346 -31
rect 373 110 390 124
rect 373 68 390 93
rect 454 122 471 139
rect 454 88 471 105
rect 498 143 515 160
rect 498 109 515 126
rect 498 71 515 92
rect 373 63 475 68
rect 498 64 532 71
rect 373 46 454 63
rect 471 46 479 63
rect 498 47 507 64
rect 524 47 532 64
rect 373 43 475 46
rect 373 20 390 43
rect 373 -14 390 3
rect 373 -39 390 -31
rect 407 -20 426 43
rect 498 41 532 47
rect 454 17 471 26
rect 407 -27 435 -20
rect 304 -57 312 -40
rect 407 -44 415 -27
rect 432 -44 435 -27
rect 407 -51 435 -44
rect 271 -58 312 -57
rect 454 -52 471 0
rect 498 17 515 41
rect 498 -10 515 0
rect 490 -36 553 -32
rect 454 -76 472 -52
rect 490 -53 495 -36
rect 512 -53 553 -36
rect 490 -57 553 -53
rect 427 -77 472 -76
rect 421 -78 472 -77
rect -144 -91 553 -78
rect -144 -108 -110 -91
rect -93 -108 -26 -91
rect -9 -108 58 -91
rect 75 -108 142 -91
rect 159 -108 226 -91
rect 243 -108 310 -91
rect 327 -108 394 -91
rect 411 -108 478 -91
rect 495 -108 553 -91
rect -144 -120 553 -108
<< viali >>
rect 136 198 153 214
rect 136 197 153 198
rect -106 46 -89 63
rect -56 47 -39 64
rect 6 46 23 63
rect 70 -46 87 -29
rect 355 152 372 169
rect 281 -40 302 -36
rect 507 47 524 64
rect 281 -57 287 -40
rect 287 -57 302 -40
rect 415 -44 432 -27
rect 495 -53 512 -36
<< metal1 >>
rect 128 218 161 221
rect 128 192 131 218
rect 158 192 161 218
rect 128 189 161 192
rect 341 169 382 182
rect -112 168 -83 169
rect 341 168 355 169
rect -113 152 355 168
rect 372 152 382 169
rect -113 136 382 152
rect -112 63 -83 136
rect -112 46 -106 63
rect -89 46 -83 63
rect -112 -29 -83 46
rect -64 70 -29 74
rect -64 44 -59 70
rect -33 44 -29 70
rect -64 39 -29 44
rect 0 64 532 69
rect 0 63 507 64
rect 0 46 6 63
rect 23 47 507 63
rect 524 47 532 64
rect 23 46 532 47
rect 0 41 532 46
rect 59 -29 98 -21
rect -112 -46 70 -29
rect 87 -46 98 -29
rect 409 -27 518 -20
rect -112 -72 98 -46
rect 275 -33 308 -30
rect 275 -60 279 -33
rect 305 -60 308 -33
rect 409 -44 415 -27
rect 432 -36 518 -27
rect 432 -44 495 -36
rect 409 -50 495 -44
rect 416 -51 495 -50
rect 490 -53 495 -51
rect 512 -53 518 -36
rect 490 -59 518 -53
rect 275 -61 308 -60
rect 276 -62 308 -61
<< via1 >>
rect 131 214 158 218
rect 131 197 136 214
rect 136 197 153 214
rect 153 197 158 214
rect 131 192 158 197
rect -59 64 -33 70
rect -59 47 -56 64
rect -56 47 -39 64
rect -39 47 -33 64
rect -59 44 -33 47
rect 279 -36 305 -33
rect 279 -57 281 -36
rect 281 -57 302 -36
rect 302 -57 305 -36
rect 279 -60 305 -57
<< metal2 >>
rect -63 218 305 221
rect -63 192 131 218
rect 158 192 305 218
rect -63 191 305 192
rect -63 74 -30 191
rect 129 189 158 191
rect -64 70 -29 74
rect -64 44 -59 70
rect -33 44 -29 70
rect -64 39 -29 44
rect 272 -28 305 191
rect 274 -33 311 -28
rect 274 -60 279 -33
rect 305 -60 311 -33
rect 274 -64 311 -60
<< labels >>
rlabel locali -144 46 -144 63 3 Clk_In
port 2 e
rlabel space -144 -121 -144 -78 3 GND
port 3 e
rlabel locali 553 -57 553 -32 7 Clk_Out
port 4 w
rlabel locali -146 236 -146 284 3 VDD
port 5 e
<< end >>
