* SPICE3 file created from PD_new.ext - technology: sky130A
.include sky130nm.lib
.option scale=0.01u

XM1000 Clk_Ref Clk_Ref a_0_161# VDD sky130_fd_pr__pfet_01v8 w=65 l=15
+  ad=2145 pd=196 as=2145 ps=196
XM1001 Up a_272_265# VDD VDD sky130_fd_pr__pfet_01v8 w=96 l=15
+  ad=2880 pd=252 as=2064.84 ps=173.327
XM1002 GND a_0_161# a_272_265# GND sky130_fd_pr__nfet_01v8 w=36 l=15
+  ad=842.4 pd=91.8 as=1116 ps=134
XM1003 a_0_105# Clk_Ref a_0_48# GND sky130_fd_pr__nfet_01v8 w=180 l=15
+  ad=4508.18 pd=301.364 as=5220 ps=370
XM1004 a_179_n156# Clk2 a_123_n156# GND sky130_fd_pr__nfet_01v8 w=84 l=15
+  ad=2772 pd=234 as=2103.82 ps=140.636
XM1005 a_315_n149# Clk2 a_123_n156# VDD sky130_fd_pr__pfet_01v8 w=65 l=15
+  ad=2145 pd=196 as=2145 ps=196
XM1006 VDD a_0_161# a_272_265# VDD sky130_fd_pr__pfet_01v8 w=72 l=15
+  ad=1548.63 pd=129.995 as=2232 ps=206
XM1007 Down a_400_n165# GND GND sky130_fd_pr__nfet_01v8 w=48 l=15
+  ad=1392 pd=154 as=1123.2 ps=122.4
XM1008 VDD Clk_Ref a_0_105# VDD sky130_fd_pr__pfet_01v8 w=65 l=15
+  ad=1398.07 pd=117.357 as=2145 ps=196
XM1009 GND a_179_n156# a_400_n165# GND sky130_fd_pr__nfet_01v8 w=36 l=15
+  ad=842.4 pd=91.8 as=1116 ps=134
XM1010 Clk2 Clk2 a_179_n156# VDD sky130_fd_pr__pfet_01v8 w=65 l=15
+  ad=2145 pd=196 as=2145 ps=196
XM1011 VDD a_179_n156# a_400_n165# VDD sky130_fd_pr__pfet_01v8 w=72 l=15
+  ad=1548.63 pd=129.995 as=2232 ps=206
XM1012 a_66_n156# Clk_Ref GND GND sky130_fd_pr__nfet_01v8 w=36 l=15
+  ad=1044 pd=74 as=842.4 ps=91.8
XM1013 Down a_400_n165# VDD VDD sky130_fd_pr__pfet_01v8 w=96 l=15
+  ad=2880 pd=252 as=2064.84 ps=173.327
XM1014 Up a_272_265# GND GND sky130_fd_pr__nfet_01v8 w=48 l=15
+  ad=1392 pd=154 as=1123.2 ps=122.4
xM1015 a_0_48# Clk2 GND GND sky130_fd_pr__nfet_01v8 w=36 l=15
+  ad=1044 pd=74 as=842.4 ps=91.8
XM1016 a_123_n156# Clk2 a_66_n156# GND sky130_fd_pr__nfet_01v8 w=180 l=15
+  ad=4508.18 pd=301.364 as=5220 ps=370
XM1017 a_0_161# Clk_Ref a_0_105# GND sky130_fd_pr__nfet_01v8 w=84 l=15
+  ad=2772 pd=234 as=2103.82 ps=140.636
C0 VDD GND 3.20fF

v1 VDD GND 1.8
v2 Clk_Ref 0 PULSE 0 1.8 40n 6p 6p 100n 200n
v3 Clk2 0 PULSE 0 1.8 6p 6p 100n 200n

.control
tran 1n 5u
plot v(Clk_Ref) v(Clk2) v(Up)+2 v(Down)+2
.endc
