*PD_10T
.include sky130nm.lib

xm1 1 clk1 3 1 sky130_fd_pr__pfet_01v8 l=150n w=420n 
xm2 3 clk1 4 0 sky130_fd_pr__nfet_01v8 l=150n w=420n
xm3 4 clk2 0 0 sky130_fd_pr__nfet_01v8 l=150n w=420n

xm4 1 clk2 6 1 sky130_fd_pr__pfet_01v8 l=150n w=420n 
xm5 6 clk2 7 0 sky130_fd_pr__nfet_01v8 l=150n w=420n
xm6 7 clk1 0 0 sky130_fd_pr__nfet_01v8 l=150n w=420n

xm7 up clk1 3 0 sky130_fd_pr__nfet_01v8 l=150n w=1440n 
xm8 clk1 clk1 up 1 sky130_fd_pr__pfet_01v8 l=150n w=1440n

xm9 down clk2 6 0 sky130_fd_pr__nfet_01v8 l=150n w=1440n
xm10 clk2 clk2 down 1 sky130_fd_pr__pfet_01v8 l=150n w=1440n


*output cap
c1 up 0 0.8f
c2 down 0 0.8f

*sources
v1 1 0 1.8v
v2 clk1 0 pulse(0 1.8 0 2ns 2ns 100ns 200ns)
v3 clk2 0 pulse(0 1.8 16ns 2ns 2ns 100ns 200ns) 

*simulation
.control
tran 10ns 800ns 120ns
plot v(clk2)+4 v(clk1)+4 v(up)+2 v(down)
.endc
.end
