magic
tech sky130A
magscale 1 2
timestamp 1607727576
<< metal1 >>
rect -1850 18798 -1474 18824
rect -1850 18744 -1812 18798
rect -1853 18513 -1812 18744
rect -1850 18456 -1812 18513
rect -1508 18744 -1474 18798
rect -1508 18513 8156 18744
rect -1508 18456 -1474 18513
rect -1850 18424 -1474 18456
rect -2846 18254 -2470 18280
rect -2846 17912 -2808 18254
rect -2504 18206 -2470 18254
rect -2504 17968 8148 18206
rect -2504 17912 -2470 17968
rect -2846 17880 -2470 17912
rect -1848 17432 -1472 17458
rect -1848 17385 -1810 17432
rect -1849 17150 -1810 17385
rect -1848 17090 -1810 17150
rect -1506 17385 -1472 17432
rect -1506 17150 8136 17385
rect -1506 17090 -1472 17150
rect -1848 17058 -1472 17090
rect -2812 16304 -2436 16330
rect -2812 15962 -2774 16304
rect -2470 16260 -2436 16304
rect -2470 16022 8132 16260
rect -2470 15962 -2436 16022
rect -2812 15930 -2436 15962
rect -1886 15180 -1510 15206
rect -1886 14838 -1848 15180
rect -1544 15134 -1510 15180
rect -1544 14896 8140 15134
rect -1544 14838 -1510 14896
rect -1886 14806 -1510 14838
rect -2846 8302 -2470 8328
rect -2846 7960 -2808 8302
rect -2504 7960 -2470 8302
rect -2846 7928 -2470 7960
<< via1 >>
rect -1812 18456 -1508 18798
rect -2808 17912 -2504 18254
rect -1810 17090 -1506 17432
rect -2774 15962 -2470 16304
rect -1848 14838 -1544 15180
rect -2808 7960 -2504 8302
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 23686 696778 23865 696780
rect 23654 696744 23900 696778
rect 23654 696742 23804 696744
rect 23654 696686 23694 696742
rect 23750 696688 23804 696742
rect 23860 696688 23900 696744
rect 23750 696686 23900 696688
rect 23654 696624 23900 696686
rect 23654 696568 23694 696624
rect 23750 696568 23804 696624
rect 23860 696568 23900 696624
rect 23654 696538 23900 696568
rect 56754 696550 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 56726 696548 56905 696550
rect 22593 639248 22836 639253
rect 22590 639214 22836 639248
rect 22590 639212 22740 639214
rect 22590 639156 22630 639212
rect 22686 639158 22740 639212
rect 22796 639158 22836 639214
rect 22686 639156 22836 639158
rect 22590 639094 22836 639156
rect 22590 639038 22630 639094
rect 22686 639038 22740 639094
rect 22796 639038 22836 639094
rect 22590 639008 22836 639038
rect 22593 611073 22836 639008
rect 23692 613556 23865 696538
rect 56694 696514 56940 696548
rect 56694 696512 56844 696514
rect 56694 696456 56734 696512
rect 56790 696458 56844 696512
rect 56900 696458 56940 696514
rect 56790 696456 56940 696458
rect 56694 696394 56940 696456
rect 56694 696338 56734 696394
rect 56790 696338 56844 696394
rect 56900 696338 56940 696394
rect 56694 696308 56940 696338
rect 121614 652202 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 678994 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 219589 678994 219837 678996
rect 251426 678994 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 186466 678992 215732 678994
rect 186466 678746 215737 678992
rect 215489 675160 215737 678746
rect 219589 678746 251540 678994
rect 219589 675462 219837 678746
rect 316286 678046 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 222147 677874 316398 678046
rect 222147 677873 316394 677874
rect 222147 675949 222320 677873
rect 121487 652172 121870 652202
rect 121487 652116 121536 652172
rect 121592 652116 121636 652172
rect 121692 652116 121738 652172
rect 121794 652116 121870 652172
rect 121487 652076 121870 652116
rect 121487 652020 121534 652076
rect 121590 652020 121636 652076
rect 121692 652020 121734 652076
rect 121790 652020 121870 652076
rect 121487 651987 121870 652020
rect 381146 651044 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 678964 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 678964 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 446098 678716 474498 678964
rect 478349 678716 511070 678964
rect 474249 674128 474497 678716
rect 478349 674314 478597 678716
rect 575818 678088 575930 704960
rect 575818 677822 575926 678088
rect 480907 677649 575926 677822
rect 480907 674567 481080 677649
rect 381019 651014 381402 651044
rect 381019 650958 381068 651014
rect 381124 650958 381168 651014
rect 381224 650958 381270 651014
rect 381326 650958 381402 651014
rect 381019 650918 381402 650958
rect 381019 650862 381066 650918
rect 381122 650862 381168 650918
rect 381224 650862 381266 650918
rect 381322 650862 381402 650918
rect 381019 650829 381402 650862
rect 559280 615996 559528 615998
rect 559276 615962 559528 615996
rect 559276 615960 559430 615962
rect 559276 615904 559320 615960
rect 559376 615906 559430 615960
rect 559486 615906 559528 615962
rect 559376 615904 559528 615906
rect 559276 615842 559528 615904
rect 559276 615786 559320 615842
rect 559376 615786 559430 615842
rect 559486 615786 559528 615842
rect 559276 615756 559528 615786
rect 23692 613383 26533 613556
rect 22592 610825 27228 611073
rect 22593 606973 22836 606974
rect 22593 606725 27236 606973
rect 22593 581858 22836 606725
rect 559276 592806 559524 615756
rect 553724 592558 559524 592806
rect 554180 588458 559524 588706
rect 554897 585975 558406 586148
rect 22593 581824 22840 581858
rect 22593 581822 22744 581824
rect 22593 581766 22634 581822
rect 22690 581768 22744 581822
rect 22800 581768 22840 581824
rect 22690 581766 22840 581768
rect 22593 581704 22840 581766
rect 22593 581648 22634 581704
rect 22690 581648 22744 581704
rect 22800 581648 22840 581704
rect 22593 581618 22840 581648
rect 22593 581617 22836 581618
rect 23900 524330 24073 524332
rect 23868 524296 24114 524330
rect 23868 524294 24018 524296
rect 23868 524238 23908 524294
rect 23964 524240 24018 524294
rect 24074 524240 24114 524296
rect 23964 524238 24114 524240
rect 23868 524176 24114 524238
rect 23868 524120 23908 524176
rect 23964 524120 24018 524176
rect 24074 524120 24114 524176
rect 23868 524090 24114 524120
rect 22590 466904 22838 466942
rect 22590 466902 22740 466904
rect 22590 466846 22630 466902
rect 22686 466848 22740 466902
rect 22796 466848 22838 466904
rect 22686 466846 22838 466848
rect 22590 466784 22838 466846
rect 22590 466728 22630 466784
rect 22686 466728 22740 466784
rect 22796 466728 22838 466784
rect 22590 439377 22838 466728
rect 23900 441860 24073 524090
rect 558233 522156 558406 585975
rect 559276 569046 559524 588458
rect 559276 569044 559426 569046
rect 559276 568988 559316 569044
rect 559372 568990 559426 569044
rect 559482 568990 559524 569046
rect 559372 568988 559524 568990
rect 559276 568926 559524 568988
rect 559276 568870 559316 568926
rect 559372 568870 559426 568926
rect 559482 568870 559524 568926
rect 559276 568828 559524 568870
rect 558192 522120 558440 522156
rect 558192 522118 558342 522120
rect 558192 522062 558232 522118
rect 558288 522064 558342 522118
rect 558398 522064 558440 522120
rect 558288 522062 558440 522064
rect 558192 522000 558440 522062
rect 558192 521944 558232 522000
rect 558288 521944 558342 522000
rect 558398 521944 558440 522000
rect 558192 521914 558440 521944
rect 558233 521886 558406 521914
rect 23900 441687 26656 441860
rect 22590 439129 27202 439377
rect 22590 435277 22838 435278
rect 22590 435029 27026 435277
rect 22590 409378 22838 435029
rect 22590 409376 22740 409378
rect 22590 409320 22630 409376
rect 22686 409322 22740 409376
rect 22796 409322 22838 409378
rect 22686 409320 22838 409322
rect 22590 409258 22838 409320
rect 22590 409202 22630 409258
rect 22686 409202 22740 409258
rect 22796 409202 22838 409258
rect 22590 409172 22838 409202
rect 559326 428280 559574 428324
rect 559326 428278 559476 428280
rect 559326 428222 559366 428278
rect 559422 428224 559476 428278
rect 559532 428224 559574 428280
rect 559422 428222 559574 428224
rect 559326 428160 559574 428222
rect 559326 428104 559366 428160
rect 559422 428104 559476 428160
rect 559532 428104 559574 428160
rect 559326 408078 559574 428104
rect 553514 407830 559574 408078
rect 559326 407828 559574 407830
rect 559326 403978 559574 403980
rect 554058 403730 559574 403978
rect 554492 401247 557940 401420
rect 557767 334478 557940 401247
rect 559326 381360 559574 403730
rect 559326 381358 559476 381360
rect 559326 381302 559366 381358
rect 559422 381304 559476 381358
rect 559532 381304 559574 381360
rect 559422 381302 559574 381304
rect 559326 381240 559574 381302
rect 559326 381184 559366 381240
rect 559422 381184 559476 381240
rect 559532 381184 559574 381240
rect 559326 381120 559574 381184
rect 557724 334442 557972 334478
rect 557724 334440 557874 334442
rect 557724 334384 557764 334440
rect 557820 334386 557874 334440
rect 557930 334386 557972 334442
rect 557820 334384 557972 334386
rect 557724 334322 557972 334384
rect 557724 334266 557764 334322
rect 557820 334266 557874 334322
rect 557930 334266 557972 334322
rect 557724 334236 557972 334266
rect 557767 334210 557940 334236
rect 559408 240636 559654 240714
rect 559406 240600 559654 240636
rect 559406 240598 559550 240600
rect 559406 240542 559440 240598
rect 559496 240544 559550 240598
rect 559606 240544 559654 240600
rect 559496 240542 559654 240544
rect 559406 240480 559654 240542
rect 559406 240424 559440 240480
rect 559496 240424 559550 240480
rect 559606 240424 559654 240480
rect 559406 240394 559654 240424
rect 559408 240370 559654 240394
rect 559408 217806 559656 240370
rect 552650 217558 559656 217806
rect 552578 213458 559656 213706
rect 553783 210975 558230 211148
rect 558057 146792 558230 210975
rect 559408 193724 559656 213458
rect 559408 193688 559660 193724
rect 559408 193686 559562 193688
rect 559408 193630 559452 193686
rect 559508 193632 559562 193686
rect 559618 193632 559660 193688
rect 559508 193630 559660 193632
rect 559408 193568 559660 193630
rect 559408 193512 559452 193568
rect 559508 193512 559562 193568
rect 559618 193512 559660 193568
rect 559408 193482 559660 193512
rect 559408 193436 559656 193482
rect 558018 146756 558266 146792
rect 558018 146754 558168 146756
rect 558018 146698 558058 146754
rect 558114 146700 558168 146754
rect 558224 146700 558266 146756
rect 558114 146698 558266 146700
rect 558018 146636 558266 146698
rect 558018 146580 558058 146636
rect 558114 146580 558168 146636
rect 558224 146580 558266 146636
rect 558018 146550 558266 146580
rect 558057 146502 558230 146550
rect 364 18960 8575 19198
rect -1830 18798 -1494 18814
rect -1830 18456 -1812 18798
rect -1508 18456 -1494 18798
rect -1830 18438 -1494 18456
rect -2826 18254 -2490 18270
rect -2826 17912 -2808 18254
rect -2504 17912 -2490 18254
rect -2826 17894 -2490 17912
rect -1828 17432 -1492 17448
rect -1828 17090 -1810 17432
rect -1506 17090 -1492 17432
rect -1828 17072 -1492 17090
rect -2792 16304 -2456 16320
rect -2792 15962 -2774 16304
rect -2470 15962 -2456 16304
rect -2792 15944 -2456 15962
rect -1866 15180 -1530 15196
rect -1866 14838 -1848 15180
rect -1544 14838 -1530 15180
rect -1866 14820 -1530 14838
rect -2826 8302 -2490 8318
rect -2826 7960 -2808 8302
rect -2504 7960 -2490 8302
rect -2826 7942 -2490 7960
rect 364 947 989 18960
rect 3096 17580 8968 17848
rect 3099 2896 3545 17580
rect 6028 16670 8897 16952
rect 6030 7017 6539 16670
rect 26535 16198 577945 16493
rect 26535 15853 575710 16198
rect 26533 15364 575710 15853
rect 23927 15186 575710 15364
rect 26533 14989 575710 15186
rect 26535 14671 575710 14989
rect 26541 14260 575710 14671
rect 577488 14260 577945 16198
rect 26541 14043 577945 14260
rect 22378 11049 22720 12097
rect 22378 11008 29129 11049
rect 22378 9946 27856 11008
rect 29088 9946 29129 11008
rect 22378 9907 29129 9946
rect 6030 6508 16220 7017
rect 3099 2450 11326 2896
rect 364 -880 791 947
rect 542 -960 791 -880
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 2450
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 553 -967 791 -960
rect 15922 -963 16220 6508
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 23694 696686 23750 696742
rect 23804 696688 23860 696744
rect 23694 696568 23750 696624
rect 23804 696568 23860 696624
rect 22630 639156 22686 639212
rect 22740 639158 22796 639214
rect 22630 639038 22686 639094
rect 22740 639038 22796 639094
rect 56734 696456 56790 696512
rect 56844 696458 56900 696514
rect 56734 696338 56790 696394
rect 56844 696338 56900 696394
rect 121536 652116 121592 652172
rect 121636 652116 121692 652172
rect 121738 652116 121794 652172
rect 121534 652020 121590 652076
rect 121636 652020 121692 652076
rect 121734 652020 121790 652076
rect 381068 650958 381124 651014
rect 381168 650958 381224 651014
rect 381270 650958 381326 651014
rect 381066 650862 381122 650918
rect 381168 650862 381224 650918
rect 381266 650862 381322 650918
rect 559320 615904 559376 615960
rect 559430 615906 559486 615962
rect 559320 615786 559376 615842
rect 559430 615786 559486 615842
rect 22634 581766 22690 581822
rect 22744 581768 22800 581824
rect 22634 581648 22690 581704
rect 22744 581648 22800 581704
rect 23908 524238 23964 524294
rect 24018 524240 24074 524296
rect 23908 524120 23964 524176
rect 24018 524120 24074 524176
rect 22630 466846 22686 466902
rect 22740 466848 22796 466904
rect 22630 466728 22686 466784
rect 22740 466728 22796 466784
rect 559316 568988 559372 569044
rect 559426 568990 559482 569046
rect 559316 568870 559372 568926
rect 559426 568870 559482 568926
rect 558232 522062 558288 522118
rect 558342 522064 558398 522120
rect 558232 521944 558288 522000
rect 558342 521944 558398 522000
rect 22630 409320 22686 409376
rect 22740 409322 22796 409378
rect 22630 409202 22686 409258
rect 22740 409202 22796 409258
rect 559366 428222 559422 428278
rect 559476 428224 559532 428280
rect 559366 428104 559422 428160
rect 559476 428104 559532 428160
rect 559366 381302 559422 381358
rect 559476 381304 559532 381360
rect 559366 381184 559422 381240
rect 559476 381184 559532 381240
rect 557764 334384 557820 334440
rect 557874 334386 557930 334442
rect 557764 334266 557820 334322
rect 557874 334266 557930 334322
rect 559440 240542 559496 240598
rect 559550 240544 559606 240600
rect 559440 240424 559496 240480
rect 559550 240424 559606 240480
rect 559452 193630 559508 193686
rect 559562 193632 559618 193688
rect 559452 193512 559508 193568
rect 559562 193512 559618 193568
rect 558058 146698 558114 146754
rect 558168 146700 558224 146756
rect 558058 146580 558114 146636
rect 558168 146580 558224 146636
rect -1808 18462 -1514 18790
rect -2804 17918 -2510 18246
rect -1806 17096 -1512 17424
rect -2770 15968 -2476 16296
rect -1844 14844 -1550 15172
rect -2804 7966 -2510 8294
rect 575710 14260 577488 16198
rect 27856 9946 29088 11008
<< metal3 >>
rect 583520 697900 584960 698140
rect -960 696744 23902 696780
rect -960 696742 23804 696744
rect -960 696686 23694 696742
rect 23750 696688 23804 696742
rect 23860 696688 23902 696744
rect 23750 696686 23902 696688
rect -960 696624 23902 696686
rect -960 696568 23694 696624
rect 23750 696568 23804 696624
rect 23860 696568 23902 696624
rect -960 696540 23902 696568
rect 23654 696538 23900 696540
rect 50407 696524 56940 696554
rect 50407 696522 50714 696524
rect 50407 696458 50462 696522
rect 50526 696458 50582 696522
rect 50646 696460 50714 696522
rect 50778 696514 56940 696524
rect 50778 696512 56844 696514
rect 50778 696460 56734 696512
rect 50646 696458 56734 696460
rect 50407 696456 56734 696458
rect 56790 696458 56844 696512
rect 56900 696458 56940 696514
rect 56790 696456 56940 696458
rect 50407 696406 56940 696456
rect 50407 696404 50712 696406
rect 50407 696340 50460 696404
rect 50524 696340 50580 696404
rect 50644 696342 50712 696404
rect 50776 696394 56940 696406
rect 50776 696342 56734 696394
rect 50644 696340 56734 696342
rect 50407 696338 56734 696340
rect 56790 696338 56844 696394
rect 56900 696338 56940 696394
rect 50407 696308 56940 696338
rect 583520 686204 584960 686444
rect -960 682124 480 682364
rect 583520 674508 584960 674748
rect -960 667844 480 668084
rect 530488 662876 584960 662916
rect 530488 662874 530802 662876
rect 530488 662810 530550 662874
rect 530614 662810 530670 662874
rect 530734 662812 530802 662874
rect 530866 662812 584960 662876
rect 530734 662810 584960 662812
rect 530488 662758 584960 662810
rect 530488 662756 530800 662758
rect 530488 662692 530548 662756
rect 530612 662692 530668 662756
rect 530732 662694 530800 662756
rect 530864 662694 584960 662758
rect 530732 662692 584960 662694
rect 530488 662676 584960 662692
rect 530496 662662 530906 662676
rect -960 653428 480 653668
rect 121465 652176 121891 652190
rect 121465 652112 121532 652176
rect 121596 652112 121632 652176
rect 121696 652112 121734 652176
rect 121798 652112 121891 652176
rect 121465 652080 121891 652112
rect 121465 652016 121530 652080
rect 121594 652016 121632 652080
rect 121696 652016 121730 652080
rect 121794 652016 121891 652080
rect 121465 652007 121891 652016
rect 380992 651018 381414 651090
rect 380992 650954 381064 651018
rect 381128 650954 381164 651018
rect 381228 650954 381266 651018
rect 381330 650954 381414 651018
rect 583520 650980 584960 651220
rect 380992 650922 381414 650954
rect 380992 650858 381062 650922
rect 381126 650858 381164 650922
rect 381228 650858 381262 650922
rect 381326 650858 381414 650922
rect 380992 650816 381414 650858
rect 583520 639284 584960 639524
rect -960 639214 22838 639252
rect -960 639212 22740 639214
rect -960 639156 22630 639212
rect 22686 639158 22740 639212
rect 22796 639158 22838 639214
rect 22686 639156 22838 639158
rect -960 639094 22838 639156
rect -960 639038 22630 639094
rect 22686 639038 22740 639094
rect 22796 639038 22838 639094
rect -960 639012 22838 639038
rect 22590 639010 22838 639012
rect 22590 639008 22836 639010
rect 583520 627588 584960 627828
rect -960 624732 480 624972
rect 559274 615962 584960 615996
rect 559274 615960 559430 615962
rect 559274 615904 559320 615960
rect 559376 615906 559430 615960
rect 559486 615906 584960 615962
rect 559376 615904 584960 615906
rect 559274 615842 584960 615904
rect 559274 615786 559320 615842
rect 559376 615786 559430 615842
rect 559486 615786 584960 615842
rect 559274 615756 584960 615786
rect -960 610316 480 610556
rect 583520 604060 584960 604300
rect -960 595900 480 596140
rect 583520 592364 584960 592604
rect -960 581824 22842 581860
rect -960 581822 22744 581824
rect -960 581766 22634 581822
rect 22690 581768 22744 581822
rect 22800 581768 22842 581824
rect 22690 581766 22842 581768
rect -960 581704 22842 581766
rect -960 581648 22634 581704
rect 22690 581648 22744 581704
rect 22800 581648 22842 581704
rect -960 581620 22842 581648
rect 22594 581618 22840 581620
rect 583520 580668 584960 580908
rect 559276 569076 559524 569080
rect 559252 569046 584960 569076
rect 559252 569044 559426 569046
rect 559252 568988 559316 569044
rect 559372 568990 559426 569044
rect 559482 568990 584960 569046
rect 559372 568988 584960 568990
rect 559252 568926 584960 568988
rect 559252 568870 559316 568926
rect 559372 568870 559426 568926
rect 559482 568870 584960 568926
rect 559252 568836 584960 568870
rect -960 567204 480 567444
rect 583520 557140 584960 557380
rect -960 552924 480 553164
rect 583520 545444 584960 545684
rect -960 538508 480 538748
rect 583520 533748 584960 533988
rect -960 524296 24116 524332
rect -960 524294 24018 524296
rect -960 524238 23908 524294
rect 23964 524240 24018 524294
rect 24074 524240 24116 524296
rect 23964 524238 24116 524240
rect -960 524176 24116 524238
rect -960 524120 23908 524176
rect 23964 524120 24018 524176
rect 24074 524120 24116 524176
rect -960 524092 24116 524120
rect 23868 524090 24114 524092
rect 558152 522120 584960 522156
rect 558152 522118 558342 522120
rect 558152 522062 558232 522118
rect 558288 522064 558342 522118
rect 558398 522064 584960 522120
rect 558288 522062 584960 522064
rect 558152 522000 584960 522062
rect 558152 521944 558232 522000
rect 558288 521944 558342 522000
rect 558398 521944 584960 522000
rect 558152 521916 584960 521944
rect 558192 521914 558440 521916
rect 583520 510220 584960 510460
rect -960 509812 480 510052
rect 583520 498524 584960 498764
rect -960 495396 480 495636
rect 583520 486692 584960 486932
rect -960 480980 480 481220
rect 530452 475236 530960 475244
rect 530446 475204 584960 475236
rect 530446 475202 530766 475204
rect 530446 475138 530514 475202
rect 530578 475138 530634 475202
rect 530698 475140 530766 475202
rect 530830 475140 584960 475204
rect 530698 475138 584960 475140
rect 530446 475086 584960 475138
rect 530446 475084 530764 475086
rect 530446 475020 530512 475084
rect 530576 475020 530632 475084
rect 530696 475022 530764 475084
rect 530828 475022 584960 475086
rect 530696 475020 584960 475022
rect 530446 474996 584960 475020
rect 530460 474990 530870 474996
rect -960 466904 22838 466940
rect -960 466902 22740 466904
rect -960 466846 22630 466902
rect 22686 466848 22740 466902
rect 22796 466848 22838 466904
rect 22686 466846 22838 466848
rect -960 466784 22838 466846
rect -960 466728 22630 466784
rect 22686 466728 22740 466784
rect 22796 466728 22838 466784
rect -960 466700 22838 466728
rect 22590 466698 22836 466700
rect 583520 463300 584960 463540
rect -960 452284 480 452524
rect 583520 451604 584960 451844
rect 583520 439772 584960 440012
rect -960 437868 480 438108
rect 559190 428280 584960 428316
rect 559190 428278 559476 428280
rect 559190 428222 559366 428278
rect 559422 428224 559476 428278
rect 559532 428224 584960 428280
rect 559422 428222 584960 428224
rect 559190 428160 584960 428222
rect 559190 428104 559366 428160
rect 559422 428104 559476 428160
rect 559532 428104 584960 428160
rect 559190 428076 584960 428104
rect 559326 428074 559574 428076
rect -960 423588 480 423828
rect 583520 416380 584960 416620
rect -960 409378 22838 409412
rect -960 409376 22740 409378
rect -960 409320 22630 409376
rect 22686 409322 22740 409376
rect 22796 409322 22838 409378
rect 22686 409320 22838 409322
rect -960 409258 22838 409320
rect -960 409202 22630 409258
rect 22686 409202 22740 409258
rect 22796 409202 22838 409258
rect -960 409172 22838 409202
rect 583520 404684 584960 404924
rect -960 394892 480 395132
rect 583520 392852 584960 393092
rect 559236 381360 584960 381396
rect 559236 381358 559476 381360
rect 559236 381302 559366 381358
rect 559422 381304 559476 381358
rect 559532 381304 584960 381360
rect 559422 381302 584960 381304
rect 559236 381240 584960 381302
rect 559236 381184 559366 381240
rect 559422 381184 559476 381240
rect 559532 381184 584960 381240
rect 559236 381156 584960 381184
rect 559326 381154 559574 381156
rect -960 380476 480 380716
rect 583520 369460 584960 369700
rect -960 366060 480 366300
rect 583520 357764 584960 358004
rect -960 351994 50322 352020
rect -960 351992 50218 351994
rect -960 351928 49966 351992
rect 50030 351928 50086 351992
rect 50150 351930 50218 351992
rect 50282 351930 50322 351994
rect 50150 351928 50322 351930
rect -960 351876 50322 351928
rect -960 351874 50216 351876
rect -960 351810 49964 351874
rect 50028 351810 50084 351874
rect 50148 351812 50216 351874
rect 50280 351812 50322 351876
rect 50148 351810 50322 351812
rect -960 351780 50322 351810
rect 583520 345932 584960 346172
rect -960 337364 480 337604
rect 557700 334442 584960 334476
rect 557700 334440 557874 334442
rect 557700 334384 557764 334440
rect 557820 334386 557874 334440
rect 557930 334386 584960 334442
rect 557820 334384 584960 334386
rect 557700 334322 584960 334384
rect 557700 334266 557764 334322
rect 557820 334266 557874 334322
rect 557930 334266 584960 334322
rect 557700 334236 584960 334266
rect -960 322948 480 323188
rect 583520 322540 584960 322780
rect 583520 310708 584960 310948
rect -960 308668 480 308908
rect 583520 299012 584960 299252
rect -960 294252 480 294492
rect 529314 287556 529772 287558
rect 529276 287518 584960 287556
rect 529276 287516 529628 287518
rect 529276 287452 529376 287516
rect 529440 287452 529496 287516
rect 529560 287454 529628 287516
rect 529692 287454 584960 287518
rect 529560 287452 584960 287454
rect 529276 287400 584960 287452
rect 529276 287398 529626 287400
rect 529276 287334 529374 287398
rect 529438 287334 529494 287398
rect 529558 287336 529626 287398
rect 529690 287336 584960 287400
rect 529558 287334 584960 287336
rect 529276 287316 584960 287334
rect 529322 287304 529732 287316
rect -960 279972 480 280212
rect 583520 275620 584960 275860
rect -960 265556 480 265796
rect 583520 263788 584960 264028
rect 583520 252092 584960 252332
rect -960 251140 480 251380
rect 559356 240600 584960 240636
rect 559356 240598 559550 240600
rect 559356 240542 559440 240598
rect 559496 240544 559550 240598
rect 559606 240544 584960 240600
rect 559496 240542 584960 240544
rect 559356 240480 584960 240542
rect 559356 240424 559440 240480
rect 559496 240424 559550 240480
rect 559606 240424 584960 240480
rect 559356 240396 584960 240424
rect 559406 240394 559654 240396
rect -960 236860 480 237100
rect 583520 228700 584960 228940
rect -960 222444 480 222684
rect 583520 216868 584960 217108
rect -960 208028 480 208268
rect 583520 205172 584960 205412
rect -960 193748 480 193988
rect 559412 193716 559660 193722
rect 559384 193688 584960 193716
rect 559384 193686 559562 193688
rect 559384 193630 559452 193686
rect 559508 193632 559562 193686
rect 559618 193632 584960 193688
rect 559508 193630 584960 193632
rect 559384 193568 584960 193630
rect 559384 193512 559452 193568
rect 559508 193512 559562 193568
rect 559618 193512 584960 193568
rect 559384 193476 584960 193512
rect 583520 181780 584960 182020
rect -960 179332 480 179572
rect 583520 169948 584960 170188
rect -960 164916 480 165156
rect 583520 158252 584960 158492
rect -960 150636 480 150876
rect 558002 146756 584960 146796
rect 558002 146754 558168 146756
rect 558002 146698 558058 146754
rect 558114 146700 558168 146754
rect 558224 146700 584960 146756
rect 558114 146698 584960 146700
rect 558002 146636 584960 146698
rect 558002 146580 558058 146636
rect 558114 146580 558168 146636
rect 558224 146580 584960 146636
rect 558002 146556 584960 146580
rect 558018 146550 558266 146556
rect -960 136220 480 136460
rect 583520 134724 584960 134964
rect 583520 123028 584960 123268
rect -960 121940 480 122180
rect 583520 111332 584960 111572
rect -960 107524 480 107764
rect 583516 99636 584960 99876
rect -960 93108 480 93348
rect 583520 87804 584960 88044
rect -960 78828 480 79068
rect 583520 76108 584960 76348
rect -960 64412 480 64652
rect 583520 64412 584960 64652
rect 583516 52716 584960 52956
rect -960 49996 480 50236
rect 583520 40884 584960 41124
rect -960 35716 480 35956
rect 583520 29188 584960 29428
rect -944 21540 29139 21758
rect -960 21300 29139 21540
rect -843 20991 29139 21300
rect -1842 18800 -1484 18820
rect -1842 18448 -1814 18800
rect -1506 18448 -1484 18800
rect -1842 18426 -1484 18448
rect -2838 18256 -2480 18276
rect -2838 17904 -2810 18256
rect -2502 17904 -2480 18256
rect -2838 17882 -2480 17904
rect -1840 17434 -1482 17454
rect -1840 17082 -1812 17434
rect -1504 17082 -1482 17434
rect -1840 17060 -1482 17082
rect -2804 16306 -2446 16326
rect -2804 15954 -2776 16306
rect -2468 15954 -2446 16306
rect -2804 15932 -2446 15954
rect -1878 15182 -1520 15202
rect -1878 14830 -1850 15182
rect -1542 14830 -1520 15182
rect -1878 14808 -1520 14830
rect 27824 11008 29139 20991
rect 583520 17492 584960 17732
rect 27824 9946 27856 11008
rect 29088 9946 29139 11008
rect 27824 9905 29139 9946
rect 575558 16318 577640 16416
rect 575558 16198 577672 16318
rect 575558 14260 575710 16198
rect 577488 14260 577672 16198
rect -2838 8304 1762 8344
rect -2838 7952 -2810 8304
rect -2502 7952 1762 8304
rect -2838 7890 1762 7952
rect 1522 7260 1762 7890
rect -960 7020 1762 7260
rect 575558 6440 577672 14260
rect 575516 5438 584984 6440
<< via3 >>
rect 50462 696458 50526 696522
rect 50582 696458 50646 696522
rect 50714 696460 50778 696524
rect 50460 696340 50524 696404
rect 50580 696340 50644 696404
rect 50712 696342 50776 696406
rect 530550 662810 530614 662874
rect 530670 662810 530734 662874
rect 530802 662812 530866 662876
rect 530548 662692 530612 662756
rect 530668 662692 530732 662756
rect 530800 662694 530864 662758
rect 121532 652172 121596 652176
rect 121532 652116 121536 652172
rect 121536 652116 121592 652172
rect 121592 652116 121596 652172
rect 121532 652112 121596 652116
rect 121632 652172 121696 652176
rect 121632 652116 121636 652172
rect 121636 652116 121692 652172
rect 121692 652116 121696 652172
rect 121632 652112 121696 652116
rect 121734 652172 121798 652176
rect 121734 652116 121738 652172
rect 121738 652116 121794 652172
rect 121794 652116 121798 652172
rect 121734 652112 121798 652116
rect 121530 652076 121594 652080
rect 121530 652020 121534 652076
rect 121534 652020 121590 652076
rect 121590 652020 121594 652076
rect 121530 652016 121594 652020
rect 121632 652076 121696 652080
rect 121632 652020 121636 652076
rect 121636 652020 121692 652076
rect 121692 652020 121696 652076
rect 121632 652016 121696 652020
rect 121730 652076 121794 652080
rect 121730 652020 121734 652076
rect 121734 652020 121790 652076
rect 121790 652020 121794 652076
rect 121730 652016 121794 652020
rect 381064 651014 381128 651018
rect 381064 650958 381068 651014
rect 381068 650958 381124 651014
rect 381124 650958 381128 651014
rect 381064 650954 381128 650958
rect 381164 651014 381228 651018
rect 381164 650958 381168 651014
rect 381168 650958 381224 651014
rect 381224 650958 381228 651014
rect 381164 650954 381228 650958
rect 381266 651014 381330 651018
rect 381266 650958 381270 651014
rect 381270 650958 381326 651014
rect 381326 650958 381330 651014
rect 381266 650954 381330 650958
rect 381062 650918 381126 650922
rect 381062 650862 381066 650918
rect 381066 650862 381122 650918
rect 381122 650862 381126 650918
rect 381062 650858 381126 650862
rect 381164 650918 381228 650922
rect 381164 650862 381168 650918
rect 381168 650862 381224 650918
rect 381224 650862 381228 650918
rect 381164 650858 381228 650862
rect 381262 650918 381326 650922
rect 381262 650862 381266 650918
rect 381266 650862 381322 650918
rect 381322 650862 381326 650918
rect 381262 650858 381326 650862
rect 530514 475138 530578 475202
rect 530634 475138 530698 475202
rect 530766 475140 530830 475204
rect 530512 475020 530576 475084
rect 530632 475020 530696 475084
rect 530764 475022 530828 475086
rect 49966 351928 50030 351992
rect 50086 351928 50150 351992
rect 50218 351930 50282 351994
rect 49964 351810 50028 351874
rect 50084 351810 50148 351874
rect 50216 351812 50280 351876
rect 529376 287452 529440 287516
rect 529496 287452 529560 287516
rect 529628 287454 529692 287518
rect 529374 287334 529438 287398
rect 529494 287334 529558 287398
rect 529626 287336 529690 287400
rect -1814 18790 -1506 18800
rect -1814 18462 -1808 18790
rect -1808 18462 -1514 18790
rect -1514 18462 -1506 18790
rect -1814 18448 -1506 18462
rect -2810 18246 -2502 18256
rect -2810 17918 -2804 18246
rect -2804 17918 -2510 18246
rect -2510 17918 -2502 18246
rect -2810 17904 -2502 17918
rect -1812 17424 -1504 17434
rect -1812 17096 -1806 17424
rect -1806 17096 -1512 17424
rect -1512 17096 -1504 17424
rect -1812 17082 -1504 17096
rect -2776 16296 -2468 16306
rect -2776 15968 -2770 16296
rect -2770 15968 -2476 16296
rect -2476 15968 -2468 16296
rect -2776 15954 -2468 15968
rect -1850 15172 -1542 15182
rect -1850 14844 -1844 15172
rect -1844 14844 -1550 15172
rect -1550 14844 -1542 15172
rect -1850 14830 -1542 14844
rect -2810 8294 -2502 8304
rect -2810 7966 -2804 8294
rect -2804 7966 -2510 8294
rect -2510 7966 -2502 8294
rect -2810 7952 -2502 7966
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 679254 -7976 710862
rect -8576 679018 -8394 679254
rect -8158 679018 -7976 679254
rect -8576 678934 -7976 679018
rect -8576 678698 -8394 678934
rect -8158 678698 -7976 678934
rect -8576 643254 -7976 678698
rect -8576 643018 -8394 643254
rect -8158 643018 -7976 643254
rect -8576 642934 -7976 643018
rect -8576 642698 -8394 642934
rect -8158 642698 -7976 642934
rect -8576 607254 -7976 642698
rect -8576 607018 -8394 607254
rect -8158 607018 -7976 607254
rect -8576 606934 -7976 607018
rect -8576 606698 -8394 606934
rect -8158 606698 -7976 606934
rect -8576 571254 -7976 606698
rect -8576 571018 -8394 571254
rect -8158 571018 -7976 571254
rect -8576 570934 -7976 571018
rect -8576 570698 -8394 570934
rect -8158 570698 -7976 570934
rect -8576 535254 -7976 570698
rect -8576 535018 -8394 535254
rect -8158 535018 -7976 535254
rect -8576 534934 -7976 535018
rect -8576 534698 -8394 534934
rect -8158 534698 -7976 534934
rect -8576 499254 -7976 534698
rect -8576 499018 -8394 499254
rect -8158 499018 -7976 499254
rect -8576 498934 -7976 499018
rect -8576 498698 -8394 498934
rect -8158 498698 -7976 498934
rect -8576 463254 -7976 498698
rect -8576 463018 -8394 463254
rect -8158 463018 -7976 463254
rect -8576 462934 -7976 463018
rect -8576 462698 -8394 462934
rect -8158 462698 -7976 462934
rect -8576 427254 -7976 462698
rect -8576 427018 -8394 427254
rect -8158 427018 -7976 427254
rect -8576 426934 -7976 427018
rect -8576 426698 -8394 426934
rect -8158 426698 -7976 426934
rect -8576 391254 -7976 426698
rect -8576 391018 -8394 391254
rect -8158 391018 -7976 391254
rect -8576 390934 -7976 391018
rect -8576 390698 -8394 390934
rect -8158 390698 -7976 390934
rect -8576 355254 -7976 390698
rect -8576 355018 -8394 355254
rect -8158 355018 -7976 355254
rect -8576 354934 -7976 355018
rect -8576 354698 -8394 354934
rect -8158 354698 -7976 354934
rect -8576 319254 -7976 354698
rect -8576 319018 -8394 319254
rect -8158 319018 -7976 319254
rect -8576 318934 -7976 319018
rect -8576 318698 -8394 318934
rect -8158 318698 -7976 318934
rect -8576 283254 -7976 318698
rect -8576 283018 -8394 283254
rect -8158 283018 -7976 283254
rect -8576 282934 -7976 283018
rect -8576 282698 -8394 282934
rect -8158 282698 -7976 282934
rect -8576 247254 -7976 282698
rect -8576 247018 -8394 247254
rect -8158 247018 -7976 247254
rect -8576 246934 -7976 247018
rect -8576 246698 -8394 246934
rect -8158 246698 -7976 246934
rect -8576 211254 -7976 246698
rect -8576 211018 -8394 211254
rect -8158 211018 -7976 211254
rect -8576 210934 -7976 211018
rect -8576 210698 -8394 210934
rect -8158 210698 -7976 210934
rect -8576 175254 -7976 210698
rect -8576 175018 -8394 175254
rect -8158 175018 -7976 175254
rect -8576 174934 -7976 175018
rect -8576 174698 -8394 174934
rect -8158 174698 -7976 174934
rect -8576 139254 -7976 174698
rect -8576 139018 -8394 139254
rect -8158 139018 -7976 139254
rect -8576 138934 -7976 139018
rect -8576 138698 -8394 138934
rect -8158 138698 -7976 138934
rect -8576 103254 -7976 138698
rect -8576 103018 -8394 103254
rect -8158 103018 -7976 103254
rect -8576 102934 -7976 103018
rect -8576 102698 -8394 102934
rect -8158 102698 -7976 102934
rect -8576 67254 -7976 102698
rect -8576 67018 -8394 67254
rect -8158 67018 -7976 67254
rect -8576 66934 -7976 67018
rect -8576 66698 -8394 66934
rect -8158 66698 -7976 66934
rect -8576 31254 -7976 66698
rect -8576 31018 -8394 31254
rect -8158 31018 -7976 31254
rect -8576 30934 -7976 31018
rect -8576 30698 -8394 30934
rect -8158 30698 -7976 30934
rect -8576 -6926 -7976 30698
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 697254 -7036 709922
rect 11604 710478 12204 711440
rect 11604 710242 11786 710478
rect 12022 710242 12204 710478
rect 11604 710158 12204 710242
rect 11604 709922 11786 710158
rect 12022 709922 12204 710158
rect -7636 697018 -7454 697254
rect -7218 697018 -7036 697254
rect -7636 696934 -7036 697018
rect -7636 696698 -7454 696934
rect -7218 696698 -7036 696934
rect -7636 661254 -7036 696698
rect -7636 661018 -7454 661254
rect -7218 661018 -7036 661254
rect -7636 660934 -7036 661018
rect -7636 660698 -7454 660934
rect -7218 660698 -7036 660934
rect -7636 625254 -7036 660698
rect -7636 625018 -7454 625254
rect -7218 625018 -7036 625254
rect -7636 624934 -7036 625018
rect -7636 624698 -7454 624934
rect -7218 624698 -7036 624934
rect -7636 589254 -7036 624698
rect -7636 589018 -7454 589254
rect -7218 589018 -7036 589254
rect -7636 588934 -7036 589018
rect -7636 588698 -7454 588934
rect -7218 588698 -7036 588934
rect -7636 553254 -7036 588698
rect -7636 553018 -7454 553254
rect -7218 553018 -7036 553254
rect -7636 552934 -7036 553018
rect -7636 552698 -7454 552934
rect -7218 552698 -7036 552934
rect -7636 517254 -7036 552698
rect -7636 517018 -7454 517254
rect -7218 517018 -7036 517254
rect -7636 516934 -7036 517018
rect -7636 516698 -7454 516934
rect -7218 516698 -7036 516934
rect -7636 481254 -7036 516698
rect -7636 481018 -7454 481254
rect -7218 481018 -7036 481254
rect -7636 480934 -7036 481018
rect -7636 480698 -7454 480934
rect -7218 480698 -7036 480934
rect -7636 445254 -7036 480698
rect -7636 445018 -7454 445254
rect -7218 445018 -7036 445254
rect -7636 444934 -7036 445018
rect -7636 444698 -7454 444934
rect -7218 444698 -7036 444934
rect -7636 409254 -7036 444698
rect -7636 409018 -7454 409254
rect -7218 409018 -7036 409254
rect -7636 408934 -7036 409018
rect -7636 408698 -7454 408934
rect -7218 408698 -7036 408934
rect -7636 373254 -7036 408698
rect -7636 373018 -7454 373254
rect -7218 373018 -7036 373254
rect -7636 372934 -7036 373018
rect -7636 372698 -7454 372934
rect -7218 372698 -7036 372934
rect -7636 337254 -7036 372698
rect -7636 337018 -7454 337254
rect -7218 337018 -7036 337254
rect -7636 336934 -7036 337018
rect -7636 336698 -7454 336934
rect -7218 336698 -7036 336934
rect -7636 301254 -7036 336698
rect -7636 301018 -7454 301254
rect -7218 301018 -7036 301254
rect -7636 300934 -7036 301018
rect -7636 300698 -7454 300934
rect -7218 300698 -7036 300934
rect -7636 265254 -7036 300698
rect -7636 265018 -7454 265254
rect -7218 265018 -7036 265254
rect -7636 264934 -7036 265018
rect -7636 264698 -7454 264934
rect -7218 264698 -7036 264934
rect -7636 229254 -7036 264698
rect -7636 229018 -7454 229254
rect -7218 229018 -7036 229254
rect -7636 228934 -7036 229018
rect -7636 228698 -7454 228934
rect -7218 228698 -7036 228934
rect -7636 193254 -7036 228698
rect -7636 193018 -7454 193254
rect -7218 193018 -7036 193254
rect -7636 192934 -7036 193018
rect -7636 192698 -7454 192934
rect -7218 192698 -7036 192934
rect -7636 157254 -7036 192698
rect -7636 157018 -7454 157254
rect -7218 157018 -7036 157254
rect -7636 156934 -7036 157018
rect -7636 156698 -7454 156934
rect -7218 156698 -7036 156934
rect -7636 121254 -7036 156698
rect -7636 121018 -7454 121254
rect -7218 121018 -7036 121254
rect -7636 120934 -7036 121018
rect -7636 120698 -7454 120934
rect -7218 120698 -7036 120934
rect -7636 85254 -7036 120698
rect -7636 85018 -7454 85254
rect -7218 85018 -7036 85254
rect -7636 84934 -7036 85018
rect -7636 84698 -7454 84934
rect -7218 84698 -7036 84934
rect -7636 49254 -7036 84698
rect -7636 49018 -7454 49254
rect -7218 49018 -7036 49254
rect -7636 48934 -7036 49018
rect -7636 48698 -7454 48934
rect -7218 48698 -7036 48934
rect -7636 13254 -7036 48698
rect -7636 13018 -7454 13254
rect -7218 13018 -7036 13254
rect -7636 12934 -7036 13018
rect -7636 12698 -7454 12934
rect -7218 12698 -7036 12934
rect -7636 -5986 -7036 12698
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 675654 -6096 708982
rect -6696 675418 -6514 675654
rect -6278 675418 -6096 675654
rect -6696 675334 -6096 675418
rect -6696 675098 -6514 675334
rect -6278 675098 -6096 675334
rect -6696 639654 -6096 675098
rect -6696 639418 -6514 639654
rect -6278 639418 -6096 639654
rect -6696 639334 -6096 639418
rect -6696 639098 -6514 639334
rect -6278 639098 -6096 639334
rect -6696 603654 -6096 639098
rect -6696 603418 -6514 603654
rect -6278 603418 -6096 603654
rect -6696 603334 -6096 603418
rect -6696 603098 -6514 603334
rect -6278 603098 -6096 603334
rect -6696 567654 -6096 603098
rect -6696 567418 -6514 567654
rect -6278 567418 -6096 567654
rect -6696 567334 -6096 567418
rect -6696 567098 -6514 567334
rect -6278 567098 -6096 567334
rect -6696 531654 -6096 567098
rect -6696 531418 -6514 531654
rect -6278 531418 -6096 531654
rect -6696 531334 -6096 531418
rect -6696 531098 -6514 531334
rect -6278 531098 -6096 531334
rect -6696 495654 -6096 531098
rect -6696 495418 -6514 495654
rect -6278 495418 -6096 495654
rect -6696 495334 -6096 495418
rect -6696 495098 -6514 495334
rect -6278 495098 -6096 495334
rect -6696 459654 -6096 495098
rect -6696 459418 -6514 459654
rect -6278 459418 -6096 459654
rect -6696 459334 -6096 459418
rect -6696 459098 -6514 459334
rect -6278 459098 -6096 459334
rect -6696 423654 -6096 459098
rect -6696 423418 -6514 423654
rect -6278 423418 -6096 423654
rect -6696 423334 -6096 423418
rect -6696 423098 -6514 423334
rect -6278 423098 -6096 423334
rect -6696 387654 -6096 423098
rect -6696 387418 -6514 387654
rect -6278 387418 -6096 387654
rect -6696 387334 -6096 387418
rect -6696 387098 -6514 387334
rect -6278 387098 -6096 387334
rect -6696 351654 -6096 387098
rect -6696 351418 -6514 351654
rect -6278 351418 -6096 351654
rect -6696 351334 -6096 351418
rect -6696 351098 -6514 351334
rect -6278 351098 -6096 351334
rect -6696 315654 -6096 351098
rect -6696 315418 -6514 315654
rect -6278 315418 -6096 315654
rect -6696 315334 -6096 315418
rect -6696 315098 -6514 315334
rect -6278 315098 -6096 315334
rect -6696 279654 -6096 315098
rect -6696 279418 -6514 279654
rect -6278 279418 -6096 279654
rect -6696 279334 -6096 279418
rect -6696 279098 -6514 279334
rect -6278 279098 -6096 279334
rect -6696 243654 -6096 279098
rect -6696 243418 -6514 243654
rect -6278 243418 -6096 243654
rect -6696 243334 -6096 243418
rect -6696 243098 -6514 243334
rect -6278 243098 -6096 243334
rect -6696 207654 -6096 243098
rect -6696 207418 -6514 207654
rect -6278 207418 -6096 207654
rect -6696 207334 -6096 207418
rect -6696 207098 -6514 207334
rect -6278 207098 -6096 207334
rect -6696 171654 -6096 207098
rect -6696 171418 -6514 171654
rect -6278 171418 -6096 171654
rect -6696 171334 -6096 171418
rect -6696 171098 -6514 171334
rect -6278 171098 -6096 171334
rect -6696 135654 -6096 171098
rect -6696 135418 -6514 135654
rect -6278 135418 -6096 135654
rect -6696 135334 -6096 135418
rect -6696 135098 -6514 135334
rect -6278 135098 -6096 135334
rect -6696 99654 -6096 135098
rect -6696 99418 -6514 99654
rect -6278 99418 -6096 99654
rect -6696 99334 -6096 99418
rect -6696 99098 -6514 99334
rect -6278 99098 -6096 99334
rect -6696 63654 -6096 99098
rect -6696 63418 -6514 63654
rect -6278 63418 -6096 63654
rect -6696 63334 -6096 63418
rect -6696 63098 -6514 63334
rect -6278 63098 -6096 63334
rect -6696 27654 -6096 63098
rect -6696 27418 -6514 27654
rect -6278 27418 -6096 27654
rect -6696 27334 -6096 27418
rect -6696 27098 -6514 27334
rect -6278 27098 -6096 27334
rect -6696 -5046 -6096 27098
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 693654 -5156 708042
rect 8004 708598 8604 709560
rect 8004 708362 8186 708598
rect 8422 708362 8604 708598
rect 8004 708278 8604 708362
rect 8004 708042 8186 708278
rect 8422 708042 8604 708278
rect -5756 693418 -5574 693654
rect -5338 693418 -5156 693654
rect -5756 693334 -5156 693418
rect -5756 693098 -5574 693334
rect -5338 693098 -5156 693334
rect -5756 657654 -5156 693098
rect -5756 657418 -5574 657654
rect -5338 657418 -5156 657654
rect -5756 657334 -5156 657418
rect -5756 657098 -5574 657334
rect -5338 657098 -5156 657334
rect -5756 621654 -5156 657098
rect -5756 621418 -5574 621654
rect -5338 621418 -5156 621654
rect -5756 621334 -5156 621418
rect -5756 621098 -5574 621334
rect -5338 621098 -5156 621334
rect -5756 585654 -5156 621098
rect -5756 585418 -5574 585654
rect -5338 585418 -5156 585654
rect -5756 585334 -5156 585418
rect -5756 585098 -5574 585334
rect -5338 585098 -5156 585334
rect -5756 549654 -5156 585098
rect -5756 549418 -5574 549654
rect -5338 549418 -5156 549654
rect -5756 549334 -5156 549418
rect -5756 549098 -5574 549334
rect -5338 549098 -5156 549334
rect -5756 513654 -5156 549098
rect -5756 513418 -5574 513654
rect -5338 513418 -5156 513654
rect -5756 513334 -5156 513418
rect -5756 513098 -5574 513334
rect -5338 513098 -5156 513334
rect -5756 477654 -5156 513098
rect -5756 477418 -5574 477654
rect -5338 477418 -5156 477654
rect -5756 477334 -5156 477418
rect -5756 477098 -5574 477334
rect -5338 477098 -5156 477334
rect -5756 441654 -5156 477098
rect -5756 441418 -5574 441654
rect -5338 441418 -5156 441654
rect -5756 441334 -5156 441418
rect -5756 441098 -5574 441334
rect -5338 441098 -5156 441334
rect -5756 405654 -5156 441098
rect -5756 405418 -5574 405654
rect -5338 405418 -5156 405654
rect -5756 405334 -5156 405418
rect -5756 405098 -5574 405334
rect -5338 405098 -5156 405334
rect -5756 369654 -5156 405098
rect -5756 369418 -5574 369654
rect -5338 369418 -5156 369654
rect -5756 369334 -5156 369418
rect -5756 369098 -5574 369334
rect -5338 369098 -5156 369334
rect -5756 333654 -5156 369098
rect -5756 333418 -5574 333654
rect -5338 333418 -5156 333654
rect -5756 333334 -5156 333418
rect -5756 333098 -5574 333334
rect -5338 333098 -5156 333334
rect -5756 297654 -5156 333098
rect -5756 297418 -5574 297654
rect -5338 297418 -5156 297654
rect -5756 297334 -5156 297418
rect -5756 297098 -5574 297334
rect -5338 297098 -5156 297334
rect -5756 261654 -5156 297098
rect -5756 261418 -5574 261654
rect -5338 261418 -5156 261654
rect -5756 261334 -5156 261418
rect -5756 261098 -5574 261334
rect -5338 261098 -5156 261334
rect -5756 225654 -5156 261098
rect -5756 225418 -5574 225654
rect -5338 225418 -5156 225654
rect -5756 225334 -5156 225418
rect -5756 225098 -5574 225334
rect -5338 225098 -5156 225334
rect -5756 189654 -5156 225098
rect -5756 189418 -5574 189654
rect -5338 189418 -5156 189654
rect -5756 189334 -5156 189418
rect -5756 189098 -5574 189334
rect -5338 189098 -5156 189334
rect -5756 153654 -5156 189098
rect -5756 153418 -5574 153654
rect -5338 153418 -5156 153654
rect -5756 153334 -5156 153418
rect -5756 153098 -5574 153334
rect -5338 153098 -5156 153334
rect -5756 117654 -5156 153098
rect -5756 117418 -5574 117654
rect -5338 117418 -5156 117654
rect -5756 117334 -5156 117418
rect -5756 117098 -5574 117334
rect -5338 117098 -5156 117334
rect -5756 81654 -5156 117098
rect -5756 81418 -5574 81654
rect -5338 81418 -5156 81654
rect -5756 81334 -5156 81418
rect -5756 81098 -5574 81334
rect -5338 81098 -5156 81334
rect -5756 45654 -5156 81098
rect -5756 45418 -5574 45654
rect -5338 45418 -5156 45654
rect -5756 45334 -5156 45418
rect -5756 45098 -5574 45334
rect -5338 45098 -5156 45334
rect -5756 9654 -5156 45098
rect -5756 9418 -5574 9654
rect -5338 9418 -5156 9654
rect -5756 9334 -5156 9418
rect -5756 9098 -5574 9334
rect -5338 9098 -5156 9334
rect -5756 -4106 -5156 9098
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 672054 -4216 707102
rect -4816 671818 -4634 672054
rect -4398 671818 -4216 672054
rect -4816 671734 -4216 671818
rect -4816 671498 -4634 671734
rect -4398 671498 -4216 671734
rect -4816 636054 -4216 671498
rect -4816 635818 -4634 636054
rect -4398 635818 -4216 636054
rect -4816 635734 -4216 635818
rect -4816 635498 -4634 635734
rect -4398 635498 -4216 635734
rect -4816 600054 -4216 635498
rect -4816 599818 -4634 600054
rect -4398 599818 -4216 600054
rect -4816 599734 -4216 599818
rect -4816 599498 -4634 599734
rect -4398 599498 -4216 599734
rect -4816 564054 -4216 599498
rect -4816 563818 -4634 564054
rect -4398 563818 -4216 564054
rect -4816 563734 -4216 563818
rect -4816 563498 -4634 563734
rect -4398 563498 -4216 563734
rect -4816 528054 -4216 563498
rect -4816 527818 -4634 528054
rect -4398 527818 -4216 528054
rect -4816 527734 -4216 527818
rect -4816 527498 -4634 527734
rect -4398 527498 -4216 527734
rect -4816 492054 -4216 527498
rect -4816 491818 -4634 492054
rect -4398 491818 -4216 492054
rect -4816 491734 -4216 491818
rect -4816 491498 -4634 491734
rect -4398 491498 -4216 491734
rect -4816 456054 -4216 491498
rect -4816 455818 -4634 456054
rect -4398 455818 -4216 456054
rect -4816 455734 -4216 455818
rect -4816 455498 -4634 455734
rect -4398 455498 -4216 455734
rect -4816 420054 -4216 455498
rect -4816 419818 -4634 420054
rect -4398 419818 -4216 420054
rect -4816 419734 -4216 419818
rect -4816 419498 -4634 419734
rect -4398 419498 -4216 419734
rect -4816 384054 -4216 419498
rect -4816 383818 -4634 384054
rect -4398 383818 -4216 384054
rect -4816 383734 -4216 383818
rect -4816 383498 -4634 383734
rect -4398 383498 -4216 383734
rect -4816 348054 -4216 383498
rect -4816 347818 -4634 348054
rect -4398 347818 -4216 348054
rect -4816 347734 -4216 347818
rect -4816 347498 -4634 347734
rect -4398 347498 -4216 347734
rect -4816 312054 -4216 347498
rect -4816 311818 -4634 312054
rect -4398 311818 -4216 312054
rect -4816 311734 -4216 311818
rect -4816 311498 -4634 311734
rect -4398 311498 -4216 311734
rect -4816 276054 -4216 311498
rect -4816 275818 -4634 276054
rect -4398 275818 -4216 276054
rect -4816 275734 -4216 275818
rect -4816 275498 -4634 275734
rect -4398 275498 -4216 275734
rect -4816 240054 -4216 275498
rect -4816 239818 -4634 240054
rect -4398 239818 -4216 240054
rect -4816 239734 -4216 239818
rect -4816 239498 -4634 239734
rect -4398 239498 -4216 239734
rect -4816 204054 -4216 239498
rect -4816 203818 -4634 204054
rect -4398 203818 -4216 204054
rect -4816 203734 -4216 203818
rect -4816 203498 -4634 203734
rect -4398 203498 -4216 203734
rect -4816 168054 -4216 203498
rect -4816 167818 -4634 168054
rect -4398 167818 -4216 168054
rect -4816 167734 -4216 167818
rect -4816 167498 -4634 167734
rect -4398 167498 -4216 167734
rect -4816 132054 -4216 167498
rect -4816 131818 -4634 132054
rect -4398 131818 -4216 132054
rect -4816 131734 -4216 131818
rect -4816 131498 -4634 131734
rect -4398 131498 -4216 131734
rect -4816 96054 -4216 131498
rect -4816 95818 -4634 96054
rect -4398 95818 -4216 96054
rect -4816 95734 -4216 95818
rect -4816 95498 -4634 95734
rect -4398 95498 -4216 95734
rect -4816 60054 -4216 95498
rect -4816 59818 -4634 60054
rect -4398 59818 -4216 60054
rect -4816 59734 -4216 59818
rect -4816 59498 -4634 59734
rect -4398 59498 -4216 59734
rect -4816 24054 -4216 59498
rect -4816 23818 -4634 24054
rect -4398 23818 -4216 24054
rect -4816 23734 -4216 23818
rect -4816 23498 -4634 23734
rect -4398 23498 -4216 23734
rect -4816 -3166 -4216 23498
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 690054 -3276 706162
rect 4404 706718 5004 707680
rect 4404 706482 4586 706718
rect 4822 706482 5004 706718
rect 4404 706398 5004 706482
rect 4404 706162 4586 706398
rect 4822 706162 5004 706398
rect -3876 689818 -3694 690054
rect -3458 689818 -3276 690054
rect -3876 689734 -3276 689818
rect -3876 689498 -3694 689734
rect -3458 689498 -3276 689734
rect -3876 654054 -3276 689498
rect -3876 653818 -3694 654054
rect -3458 653818 -3276 654054
rect -3876 653734 -3276 653818
rect -3876 653498 -3694 653734
rect -3458 653498 -3276 653734
rect -3876 618054 -3276 653498
rect -3876 617818 -3694 618054
rect -3458 617818 -3276 618054
rect -3876 617734 -3276 617818
rect -3876 617498 -3694 617734
rect -3458 617498 -3276 617734
rect -3876 582054 -3276 617498
rect -3876 581818 -3694 582054
rect -3458 581818 -3276 582054
rect -3876 581734 -3276 581818
rect -3876 581498 -3694 581734
rect -3458 581498 -3276 581734
rect -3876 546054 -3276 581498
rect -3876 545818 -3694 546054
rect -3458 545818 -3276 546054
rect -3876 545734 -3276 545818
rect -3876 545498 -3694 545734
rect -3458 545498 -3276 545734
rect -3876 510054 -3276 545498
rect -3876 509818 -3694 510054
rect -3458 509818 -3276 510054
rect -3876 509734 -3276 509818
rect -3876 509498 -3694 509734
rect -3458 509498 -3276 509734
rect -3876 474054 -3276 509498
rect -3876 473818 -3694 474054
rect -3458 473818 -3276 474054
rect -3876 473734 -3276 473818
rect -3876 473498 -3694 473734
rect -3458 473498 -3276 473734
rect -3876 438054 -3276 473498
rect -3876 437818 -3694 438054
rect -3458 437818 -3276 438054
rect -3876 437734 -3276 437818
rect -3876 437498 -3694 437734
rect -3458 437498 -3276 437734
rect -3876 402054 -3276 437498
rect -3876 401818 -3694 402054
rect -3458 401818 -3276 402054
rect -3876 401734 -3276 401818
rect -3876 401498 -3694 401734
rect -3458 401498 -3276 401734
rect -3876 366054 -3276 401498
rect -3876 365818 -3694 366054
rect -3458 365818 -3276 366054
rect -3876 365734 -3276 365818
rect -3876 365498 -3694 365734
rect -3458 365498 -3276 365734
rect -3876 330054 -3276 365498
rect -3876 329818 -3694 330054
rect -3458 329818 -3276 330054
rect -3876 329734 -3276 329818
rect -3876 329498 -3694 329734
rect -3458 329498 -3276 329734
rect -3876 294054 -3276 329498
rect -3876 293818 -3694 294054
rect -3458 293818 -3276 294054
rect -3876 293734 -3276 293818
rect -3876 293498 -3694 293734
rect -3458 293498 -3276 293734
rect -3876 258054 -3276 293498
rect -3876 257818 -3694 258054
rect -3458 257818 -3276 258054
rect -3876 257734 -3276 257818
rect -3876 257498 -3694 257734
rect -3458 257498 -3276 257734
rect -3876 222054 -3276 257498
rect -3876 221818 -3694 222054
rect -3458 221818 -3276 222054
rect -3876 221734 -3276 221818
rect -3876 221498 -3694 221734
rect -3458 221498 -3276 221734
rect -3876 186054 -3276 221498
rect -3876 185818 -3694 186054
rect -3458 185818 -3276 186054
rect -3876 185734 -3276 185818
rect -3876 185498 -3694 185734
rect -3458 185498 -3276 185734
rect -3876 150054 -3276 185498
rect -3876 149818 -3694 150054
rect -3458 149818 -3276 150054
rect -3876 149734 -3276 149818
rect -3876 149498 -3694 149734
rect -3458 149498 -3276 149734
rect -3876 114054 -3276 149498
rect -3876 113818 -3694 114054
rect -3458 113818 -3276 114054
rect -3876 113734 -3276 113818
rect -3876 113498 -3694 113734
rect -3458 113498 -3276 113734
rect -3876 78054 -3276 113498
rect -3876 77818 -3694 78054
rect -3458 77818 -3276 78054
rect -3876 77734 -3276 77818
rect -3876 77498 -3694 77734
rect -3458 77498 -3276 77734
rect -3876 42054 -3276 77498
rect -3876 41818 -3694 42054
rect -3458 41818 -3276 42054
rect -3876 41734 -3276 41818
rect -3876 41498 -3694 41734
rect -3458 41498 -3276 41734
rect -3876 6054 -3276 41498
rect -3876 5818 -3694 6054
rect -3458 5818 -3276 6054
rect -3876 5734 -3276 5818
rect -3876 5498 -3694 5734
rect -3458 5498 -3276 5734
rect -3876 -2226 -3276 5498
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 18256 -2336 19898
rect -2936 17904 -2810 18256
rect -2502 17904 -2336 18256
rect -2936 16306 -2336 17904
rect -2936 15954 -2776 16306
rect -2468 15954 -2336 16306
rect -2936 8304 -2336 15954
rect -2936 7952 -2810 8304
rect -2502 7952 -2336 8304
rect -2936 -1286 -2336 7952
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 703520 1404 704282
rect 4404 703520 5004 706162
rect 8004 703520 8604 708042
rect 11604 703520 12204 709922
rect 29604 711418 30204 711440
rect 29604 711182 29786 711418
rect 30022 711182 30204 711418
rect 29604 711098 30204 711182
rect 29604 710862 29786 711098
rect 30022 710862 30204 711098
rect 26004 709538 26604 709560
rect 26004 709302 26186 709538
rect 26422 709302 26604 709538
rect 26004 709218 26604 709302
rect 26004 708982 26186 709218
rect 26422 708982 26604 709218
rect 22404 707658 23004 707680
rect 22404 707422 22586 707658
rect 22822 707422 23004 707658
rect 22404 707338 23004 707422
rect 22404 707102 22586 707338
rect 22822 707102 23004 707338
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 703520 19404 705222
rect 22404 703520 23004 707102
rect 26004 703520 26604 708982
rect 29604 703520 30204 710862
rect 47604 710478 48204 711440
rect 47604 710242 47786 710478
rect 48022 710242 48204 710478
rect 47604 710158 48204 710242
rect 47604 709922 47786 710158
rect 48022 709922 48204 710158
rect 44004 708598 44604 709560
rect 44004 708362 44186 708598
rect 44422 708362 44604 708598
rect 44004 708278 44604 708362
rect 44004 708042 44186 708278
rect 44422 708042 44604 708278
rect 40404 706718 41004 707680
rect 40404 706482 40586 706718
rect 40822 706482 41004 706718
rect 40404 706398 41004 706482
rect 40404 706162 40586 706398
rect 40822 706162 41004 706398
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect 34954 619530 35554 619532
rect 36804 619530 37404 704282
rect 40404 703520 41004 706162
rect 44004 703520 44604 708042
rect 47604 703520 48204 709922
rect 65604 711418 66204 711440
rect 65604 711182 65786 711418
rect 66022 711182 66204 711418
rect 65604 711098 66204 711182
rect 65604 710862 65786 711098
rect 66022 710862 66204 711098
rect 62004 709538 62604 709560
rect 62004 709302 62186 709538
rect 62422 709302 62604 709538
rect 62004 709218 62604 709302
rect 62004 708982 62186 709218
rect 62422 708982 62604 709218
rect 58404 707658 59004 707680
rect 58404 707422 58586 707658
rect 58822 707422 59004 707658
rect 58404 707338 59004 707422
rect 58404 707102 58586 707338
rect 58822 707102 59004 707338
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 703520 55404 705222
rect 58404 703520 59004 707102
rect 62004 703520 62604 708982
rect 65604 703520 66204 710862
rect 83604 710478 84204 711440
rect 83604 710242 83786 710478
rect 84022 710242 84204 710478
rect 83604 710158 84204 710242
rect 83604 709922 83786 710158
rect 84022 709922 84204 710158
rect 80004 708598 80604 709560
rect 80004 708362 80186 708598
rect 80422 708362 80604 708598
rect 80004 708278 80604 708362
rect 80004 708042 80186 708278
rect 80422 708042 80604 708278
rect 76404 706718 77004 707680
rect 76404 706482 76586 706718
rect 76822 706482 77004 706718
rect 76404 706398 77004 706482
rect 76404 706162 76586 706398
rect 76822 706162 77004 706398
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 703520 73404 704282
rect 76404 703520 77004 706162
rect 80004 703520 80604 708042
rect 83604 703520 84204 709922
rect 101604 711418 102204 711440
rect 101604 711182 101786 711418
rect 102022 711182 102204 711418
rect 101604 711098 102204 711182
rect 101604 710862 101786 711098
rect 102022 710862 102204 711098
rect 98004 709538 98604 709560
rect 98004 709302 98186 709538
rect 98422 709302 98604 709538
rect 98004 709218 98604 709302
rect 98004 708982 98186 709218
rect 98422 708982 98604 709218
rect 94404 707658 95004 707680
rect 94404 707422 94586 707658
rect 94822 707422 95004 707658
rect 94404 707338 95004 707422
rect 94404 707102 94586 707338
rect 94822 707102 95004 707338
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 703520 91404 705222
rect 94404 703520 95004 707102
rect 98004 703520 98604 708982
rect 101604 703520 102204 710862
rect 119604 710478 120204 711440
rect 119604 710242 119786 710478
rect 120022 710242 120204 710478
rect 119604 710158 120204 710242
rect 119604 709922 119786 710158
rect 120022 709922 120204 710158
rect 116004 708598 116604 709560
rect 116004 708362 116186 708598
rect 116422 708362 116604 708598
rect 116004 708278 116604 708362
rect 116004 708042 116186 708278
rect 116422 708042 116604 708278
rect 112404 706718 113004 707680
rect 112404 706482 112586 706718
rect 112822 706482 113004 706718
rect 112404 706398 113004 706482
rect 112404 706162 112586 706398
rect 112822 706162 113004 706398
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 703520 109404 704282
rect 112404 703520 113004 706162
rect 116004 703520 116604 708042
rect 119604 703520 120204 709922
rect 137604 711418 138204 711440
rect 137604 711182 137786 711418
rect 138022 711182 138204 711418
rect 137604 711098 138204 711182
rect 137604 710862 137786 711098
rect 138022 710862 138204 711098
rect 134004 709538 134604 709560
rect 134004 709302 134186 709538
rect 134422 709302 134604 709538
rect 134004 709218 134604 709302
rect 134004 708982 134186 709218
rect 134422 708982 134604 709218
rect 130404 707658 131004 707680
rect 130404 707422 130586 707658
rect 130822 707422 131004 707658
rect 130404 707338 131004 707422
rect 130404 707102 130586 707338
rect 130822 707102 131004 707338
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 703520 127404 705222
rect 130404 703520 131004 707102
rect 134004 703520 134604 708982
rect 137604 703520 138204 710862
rect 155604 710478 156204 711440
rect 155604 710242 155786 710478
rect 156022 710242 156204 710478
rect 155604 710158 156204 710242
rect 155604 709922 155786 710158
rect 156022 709922 156204 710158
rect 152004 708598 152604 709560
rect 152004 708362 152186 708598
rect 152422 708362 152604 708598
rect 152004 708278 152604 708362
rect 152004 708042 152186 708278
rect 152422 708042 152604 708278
rect 148404 706718 149004 707680
rect 148404 706482 148586 706718
rect 148822 706482 149004 706718
rect 148404 706398 149004 706482
rect 148404 706162 148586 706398
rect 148822 706162 149004 706398
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 703520 145404 704282
rect 148404 703520 149004 706162
rect 152004 703520 152604 708042
rect 155604 703520 156204 709922
rect 173604 711418 174204 711440
rect 173604 711182 173786 711418
rect 174022 711182 174204 711418
rect 173604 711098 174204 711182
rect 173604 710862 173786 711098
rect 174022 710862 174204 711098
rect 170004 709538 170604 709560
rect 170004 709302 170186 709538
rect 170422 709302 170604 709538
rect 170004 709218 170604 709302
rect 170004 708982 170186 709218
rect 170422 708982 170604 709218
rect 166404 707658 167004 707680
rect 166404 707422 166586 707658
rect 166822 707422 167004 707658
rect 166404 707338 167004 707422
rect 166404 707102 166586 707338
rect 166822 707102 167004 707338
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 703520 163404 705222
rect 166404 703520 167004 707102
rect 170004 703520 170604 708982
rect 173604 703520 174204 710862
rect 191604 710478 192204 711440
rect 191604 710242 191786 710478
rect 192022 710242 192204 710478
rect 191604 710158 192204 710242
rect 191604 709922 191786 710158
rect 192022 709922 192204 710158
rect 188004 708598 188604 709560
rect 188004 708362 188186 708598
rect 188422 708362 188604 708598
rect 188004 708278 188604 708362
rect 188004 708042 188186 708278
rect 188422 708042 188604 708278
rect 184404 706718 185004 707680
rect 184404 706482 184586 706718
rect 184822 706482 185004 706718
rect 184404 706398 185004 706482
rect 184404 706162 184586 706398
rect 184822 706162 185004 706398
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 703520 181404 704282
rect 184404 703520 185004 706162
rect 188004 703520 188604 708042
rect 191604 703520 192204 709922
rect 209604 711418 210204 711440
rect 209604 711182 209786 711418
rect 210022 711182 210204 711418
rect 209604 711098 210204 711182
rect 209604 710862 209786 711098
rect 210022 710862 210204 711098
rect 206004 709538 206604 709560
rect 206004 709302 206186 709538
rect 206422 709302 206604 709538
rect 206004 709218 206604 709302
rect 206004 708982 206186 709218
rect 206422 708982 206604 709218
rect 202404 707658 203004 707680
rect 202404 707422 202586 707658
rect 202822 707422 203004 707658
rect 202404 707338 203004 707422
rect 202404 707102 202586 707338
rect 202822 707102 203004 707338
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 34954 618930 37404 619530
rect 50416 696524 50816 696554
rect 50416 696522 50714 696524
rect 50416 696458 50462 696522
rect 50526 696458 50582 696522
rect 50646 696460 50714 696522
rect 50778 696460 50816 696524
rect 50646 696458 50816 696460
rect 50416 696406 50816 696458
rect 50416 696404 50712 696406
rect 50416 696340 50460 696404
rect 50524 696340 50580 696404
rect 50644 696342 50712 696404
rect 50776 696342 50816 696406
rect 50644 696340 50816 696342
rect 34954 614036 35554 618930
rect -1996 578454 -1396 613898
rect 50416 606762 50816 696340
rect 198804 667478 199404 705222
rect 202404 703520 203004 707102
rect 206004 703520 206604 708982
rect 209604 703520 210204 710862
rect 227604 710478 228204 711440
rect 227604 710242 227786 710478
rect 228022 710242 228204 710478
rect 227604 710158 228204 710242
rect 227604 709922 227786 710158
rect 228022 709922 228204 710158
rect 224004 708598 224604 709560
rect 224004 708362 224186 708598
rect 224422 708362 224604 708598
rect 224004 708278 224604 708362
rect 224004 708042 224186 708278
rect 224422 708042 224604 708278
rect 220404 706718 221004 707680
rect 220404 706482 220586 706718
rect 220822 706482 221004 706718
rect 220404 706398 221004 706482
rect 220404 706162 220586 706398
rect 220822 706162 221004 706398
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 703520 217404 704282
rect 220404 703520 221004 706162
rect 224004 703520 224604 708042
rect 227604 703520 228204 709922
rect 245604 711418 246204 711440
rect 245604 711182 245786 711418
rect 246022 711182 246204 711418
rect 245604 711098 246204 711182
rect 245604 710862 245786 711098
rect 246022 710862 246204 711098
rect 242004 709538 242604 709560
rect 242004 709302 242186 709538
rect 242422 709302 242604 709538
rect 242004 709218 242604 709302
rect 242004 708982 242186 709218
rect 242422 708982 242604 709218
rect 238404 707658 239004 707680
rect 238404 707422 238586 707658
rect 238822 707422 239004 707658
rect 238404 707338 239004 707422
rect 238404 707102 238586 707338
rect 238822 707102 239004 707338
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 703520 235404 705222
rect 238404 703520 239004 707102
rect 242004 703520 242604 708982
rect 245604 703520 246204 710862
rect 263604 710478 264204 711440
rect 263604 710242 263786 710478
rect 264022 710242 264204 710478
rect 263604 710158 264204 710242
rect 263604 709922 263786 710158
rect 264022 709922 264204 710158
rect 260004 708598 260604 709560
rect 260004 708362 260186 708598
rect 260422 708362 260604 708598
rect 260004 708278 260604 708362
rect 260004 708042 260186 708278
rect 260422 708042 260604 708278
rect 256404 706718 257004 707680
rect 256404 706482 256586 706718
rect 256822 706482 257004 706718
rect 256404 706398 257004 706482
rect 256404 706162 256586 706398
rect 256822 706162 257004 706398
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 667792 253404 704282
rect 256404 703520 257004 706162
rect 260004 703520 260604 708042
rect 263604 703520 264204 709922
rect 281604 711418 282204 711440
rect 281604 711182 281786 711418
rect 282022 711182 282204 711418
rect 281604 711098 282204 711182
rect 281604 710862 281786 711098
rect 282022 710862 282204 711098
rect 278004 709538 278604 709560
rect 278004 709302 278186 709538
rect 278422 709302 278604 709538
rect 278004 709218 278604 709302
rect 278004 708982 278186 709218
rect 278422 708982 278604 709218
rect 274404 707658 275004 707680
rect 274404 707422 274586 707658
rect 274822 707422 275004 707658
rect 274404 707338 275004 707422
rect 274404 707102 274586 707338
rect 274822 707102 275004 707338
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 703520 271404 705222
rect 274404 703520 275004 707102
rect 278004 703520 278604 708982
rect 281604 703520 282204 710862
rect 299604 710478 300204 711440
rect 299604 710242 299786 710478
rect 300022 710242 300204 710478
rect 299604 710158 300204 710242
rect 299604 709922 299786 710158
rect 300022 709922 300204 710158
rect 296004 708598 296604 709560
rect 296004 708362 296186 708598
rect 296422 708362 296604 708598
rect 296004 708278 296604 708362
rect 296004 708042 296186 708278
rect 296422 708042 296604 708278
rect 292404 706718 293004 707680
rect 292404 706482 292586 706718
rect 292822 706482 293004 706718
rect 292404 706398 293004 706482
rect 292404 706162 292586 706398
rect 292822 706162 293004 706398
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 703520 289404 704282
rect 292404 703520 293004 706162
rect 296004 703520 296604 708042
rect 299604 703520 300204 709922
rect 317604 711418 318204 711440
rect 317604 711182 317786 711418
rect 318022 711182 318204 711418
rect 317604 711098 318204 711182
rect 317604 710862 317786 711098
rect 318022 710862 318204 711098
rect 314004 709538 314604 709560
rect 314004 709302 314186 709538
rect 314422 709302 314604 709538
rect 314004 709218 314604 709302
rect 314004 708982 314186 709218
rect 314422 708982 314604 709218
rect 310404 707658 311004 707680
rect 310404 707422 310586 707658
rect 310822 707422 311004 707658
rect 310404 707338 311004 707422
rect 310404 707102 310586 707338
rect 310822 707102 311004 707338
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 703520 307404 705222
rect 310404 703520 311004 707102
rect 314004 703520 314604 708982
rect 317604 703520 318204 710862
rect 335604 710478 336204 711440
rect 335604 710242 335786 710478
rect 336022 710242 336204 710478
rect 335604 710158 336204 710242
rect 335604 709922 335786 710158
rect 336022 709922 336204 710158
rect 332004 708598 332604 709560
rect 332004 708362 332186 708598
rect 332422 708362 332604 708598
rect 332004 708278 332604 708362
rect 332004 708042 332186 708278
rect 332422 708042 332604 708278
rect 328404 706718 329004 707680
rect 328404 706482 328586 706718
rect 328822 706482 329004 706718
rect 328404 706398 329004 706482
rect 328404 706162 328586 706398
rect 328822 706162 329004 706398
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 703520 325404 704282
rect 328404 703520 329004 706162
rect 332004 703520 332604 708042
rect 335604 703520 336204 709922
rect 353604 711418 354204 711440
rect 353604 711182 353786 711418
rect 354022 711182 354204 711418
rect 353604 711098 354204 711182
rect 353604 710862 353786 711098
rect 354022 710862 354204 711098
rect 350004 709538 350604 709560
rect 350004 709302 350186 709538
rect 350422 709302 350604 709538
rect 350004 709218 350604 709302
rect 350004 708982 350186 709218
rect 350422 708982 350604 709218
rect 346404 707658 347004 707680
rect 346404 707422 346586 707658
rect 346822 707422 347004 707658
rect 346404 707338 347004 707422
rect 346404 707102 346586 707338
rect 346822 707102 347004 707338
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 703520 343404 705222
rect 346404 703520 347004 707102
rect 350004 703520 350604 708982
rect 353604 703520 354204 710862
rect 371604 710478 372204 711440
rect 371604 710242 371786 710478
rect 372022 710242 372204 710478
rect 371604 710158 372204 710242
rect 371604 709922 371786 710158
rect 372022 709922 372204 710158
rect 368004 708598 368604 709560
rect 368004 708362 368186 708598
rect 368422 708362 368604 708598
rect 368004 708278 368604 708362
rect 368004 708042 368186 708278
rect 368422 708042 368604 708278
rect 364404 706718 365004 707680
rect 364404 706482 364586 706718
rect 364822 706482 365004 706718
rect 364404 706398 365004 706482
rect 364404 706162 364586 706398
rect 364822 706162 365004 706398
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 703520 361404 704282
rect 364404 703520 365004 706162
rect 368004 703520 368604 708042
rect 371604 703520 372204 709922
rect 389604 711418 390204 711440
rect 389604 711182 389786 711418
rect 390022 711182 390204 711418
rect 389604 711098 390204 711182
rect 389604 710862 389786 711098
rect 390022 710862 390204 711098
rect 386004 709538 386604 709560
rect 386004 709302 386186 709538
rect 386422 709302 386604 709538
rect 386004 709218 386604 709302
rect 386004 708982 386186 709218
rect 386422 708982 386604 709218
rect 382404 707658 383004 707680
rect 382404 707422 382586 707658
rect 382822 707422 383004 707658
rect 382404 707338 383004 707422
rect 382404 707102 382586 707338
rect 382822 707102 383004 707338
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 703520 379404 705222
rect 382404 703520 383004 707102
rect 386004 703520 386604 708982
rect 389604 703520 390204 710862
rect 407604 710478 408204 711440
rect 407604 710242 407786 710478
rect 408022 710242 408204 710478
rect 407604 710158 408204 710242
rect 407604 709922 407786 710158
rect 408022 709922 408204 710158
rect 404004 708598 404604 709560
rect 404004 708362 404186 708598
rect 404422 708362 404604 708598
rect 404004 708278 404604 708362
rect 404004 708042 404186 708278
rect 404422 708042 404604 708278
rect 400404 706718 401004 707680
rect 400404 706482 400586 706718
rect 400822 706482 401004 706718
rect 400404 706398 401004 706482
rect 400404 706162 400586 706398
rect 400822 706162 401004 706398
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 703520 397404 704282
rect 400404 703520 401004 706162
rect 404004 703520 404604 708042
rect 407604 703520 408204 709922
rect 425604 711418 426204 711440
rect 425604 711182 425786 711418
rect 426022 711182 426204 711418
rect 425604 711098 426204 711182
rect 425604 710862 425786 711098
rect 426022 710862 426204 711098
rect 422004 709538 422604 709560
rect 422004 709302 422186 709538
rect 422422 709302 422604 709538
rect 422004 709218 422604 709302
rect 422004 708982 422186 709218
rect 422422 708982 422604 709218
rect 418404 707658 419004 707680
rect 418404 707422 418586 707658
rect 418822 707422 419004 707658
rect 418404 707338 419004 707422
rect 418404 707102 418586 707338
rect 418822 707102 419004 707338
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 703520 415404 705222
rect 418404 703520 419004 707102
rect 422004 703520 422604 708982
rect 425604 703520 426204 710862
rect 443604 710478 444204 711440
rect 443604 710242 443786 710478
rect 444022 710242 444204 710478
rect 443604 710158 444204 710242
rect 443604 709922 443786 710158
rect 444022 709922 444204 710158
rect 440004 708598 440604 709560
rect 440004 708362 440186 708598
rect 440422 708362 440604 708598
rect 440004 708278 440604 708362
rect 440004 708042 440186 708278
rect 440422 708042 440604 708278
rect 436404 706718 437004 707680
rect 436404 706482 436586 706718
rect 436822 706482 437004 706718
rect 436404 706398 437004 706482
rect 436404 706162 436586 706398
rect 436822 706162 437004 706398
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 703520 433404 704282
rect 436404 703520 437004 706162
rect 440004 703520 440604 708042
rect 443604 703520 444204 709922
rect 461604 711418 462204 711440
rect 461604 711182 461786 711418
rect 462022 711182 462204 711418
rect 461604 711098 462204 711182
rect 461604 710862 461786 711098
rect 462022 710862 462204 711098
rect 458004 709538 458604 709560
rect 458004 709302 458186 709538
rect 458422 709302 458604 709538
rect 458004 709218 458604 709302
rect 458004 708982 458186 709218
rect 458422 708982 458604 709218
rect 454404 707658 455004 707680
rect 454404 707422 454586 707658
rect 454822 707422 455004 707658
rect 454404 707338 455004 707422
rect 454404 707102 454586 707338
rect 454822 707102 455004 707338
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 198802 666878 211166 667478
rect 222664 667192 253408 667792
rect 450804 666146 451404 705222
rect 454404 703520 455004 707102
rect 458004 703520 458604 708982
rect 461604 703520 462204 710862
rect 479604 710478 480204 711440
rect 479604 710242 479786 710478
rect 480022 710242 480204 710478
rect 479604 710158 480204 710242
rect 479604 709922 479786 710158
rect 480022 709922 480204 710158
rect 476004 708598 476604 709560
rect 476004 708362 476186 708598
rect 476422 708362 476604 708598
rect 476004 708278 476604 708362
rect 476004 708042 476186 708278
rect 476422 708042 476604 708278
rect 472404 706718 473004 707680
rect 472404 706482 472586 706718
rect 472822 706482 473004 706718
rect 472404 706398 473004 706482
rect 472404 706162 472586 706398
rect 472822 706162 473004 706398
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 703520 469404 704282
rect 472404 703520 473004 706162
rect 476004 703520 476604 708042
rect 479604 703520 480204 709922
rect 497604 711418 498204 711440
rect 497604 711182 497786 711418
rect 498022 711182 498204 711418
rect 497604 711098 498204 711182
rect 497604 710862 497786 711098
rect 498022 710862 498204 711098
rect 494004 709538 494604 709560
rect 494004 709302 494186 709538
rect 494422 709302 494604 709538
rect 494004 709218 494604 709302
rect 494004 708982 494186 709218
rect 494422 708982 494604 709218
rect 490404 707658 491004 707680
rect 490404 707422 490586 707658
rect 490822 707422 491004 707658
rect 490404 707338 491004 707422
rect 490404 707102 490586 707338
rect 490822 707102 491004 707338
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 703520 487404 705222
rect 490404 703520 491004 707102
rect 494004 703520 494604 708982
rect 497604 703520 498204 710862
rect 515604 710478 516204 711440
rect 515604 710242 515786 710478
rect 516022 710242 516204 710478
rect 515604 710158 516204 710242
rect 515604 709922 515786 710158
rect 516022 709922 516204 710158
rect 512004 708598 512604 709560
rect 512004 708362 512186 708598
rect 512422 708362 512604 708598
rect 512004 708278 512604 708362
rect 512004 708042 512186 708278
rect 512422 708042 512604 708278
rect 508404 706718 509004 707680
rect 508404 706482 508586 706718
rect 508822 706482 509004 706718
rect 508404 706398 509004 706482
rect 508404 706162 508586 706398
rect 508822 706162 509004 706398
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 666616 505404 704282
rect 508404 703520 509004 706162
rect 512004 703520 512604 708042
rect 515604 703520 516204 709922
rect 533604 711418 534204 711440
rect 533604 711182 533786 711418
rect 534022 711182 534204 711418
rect 533604 711098 534204 711182
rect 533604 710862 533786 711098
rect 534022 710862 534204 711098
rect 530004 709538 530604 709560
rect 530004 709302 530186 709538
rect 530422 709302 530604 709538
rect 530004 709218 530604 709302
rect 530004 708982 530186 709218
rect 530422 708982 530604 709218
rect 526404 707658 527004 707680
rect 526404 707422 526586 707658
rect 526822 707422 527004 707658
rect 526404 707338 527004 707422
rect 526404 707102 526586 707338
rect 526822 707102 527004 707338
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 703520 523404 705222
rect 526404 703520 527004 707102
rect 530004 703520 530604 708982
rect 533604 703520 534204 710862
rect 551604 710478 552204 711440
rect 551604 710242 551786 710478
rect 552022 710242 552204 710478
rect 551604 710158 552204 710242
rect 551604 709922 551786 710158
rect 552022 709922 552204 710158
rect 548004 708598 548604 709560
rect 548004 708362 548186 708598
rect 548422 708362 548604 708598
rect 548004 708278 548604 708362
rect 548004 708042 548186 708278
rect 548422 708042 548604 708278
rect 544404 706718 545004 707680
rect 544404 706482 544586 706718
rect 544822 706482 545004 706718
rect 544404 706398 545004 706482
rect 544404 706162 544586 706398
rect 544822 706162 545004 706398
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 703520 541404 704282
rect 544404 703520 545004 706162
rect 548004 703520 548604 708042
rect 551604 703520 552204 709922
rect 569604 711418 570204 711440
rect 569604 711182 569786 711418
rect 570022 711182 570204 711418
rect 569604 711098 570204 711182
rect 569604 710862 569786 711098
rect 570022 710862 570204 711098
rect 566004 709538 566604 709560
rect 566004 709302 566186 709538
rect 566422 709302 566604 709538
rect 566004 709218 566604 709302
rect 566004 708982 566186 709218
rect 566422 708982 566604 709218
rect 562404 707658 563004 707680
rect 562404 707422 562586 707658
rect 562822 707422 563004 707658
rect 562404 707338 563004 707422
rect 562404 707102 562586 707338
rect 562822 707102 563004 707338
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 703520 559404 705222
rect 562404 703520 563004 707102
rect 566004 703520 566604 708982
rect 569604 703520 570204 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect 580404 706718 581004 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 580404 706482 580586 706718
rect 580822 706482 581004 706718
rect 580404 706398 581004 706482
rect 580404 706162 580586 706398
rect 580822 706162 581004 706398
rect 576804 704838 577404 705800
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 703520 577404 704282
rect 580404 703520 581004 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 450804 665546 469618 666146
rect 481606 666016 505410 666616
rect 450804 665540 451404 665546
rect 530510 662906 530910 662926
rect 530506 662876 530910 662906
rect 530506 662874 530802 662876
rect 530506 662810 530550 662874
rect 530614 662810 530670 662874
rect 530734 662812 530802 662874
rect 530866 662812 530910 662876
rect 530734 662810 530910 662812
rect 530506 662758 530910 662810
rect 530506 662756 530800 662758
rect 530506 662692 530548 662756
rect 530612 662692 530668 662756
rect 530732 662694 530800 662756
rect 530864 662694 530910 662758
rect 530732 662692 530910 662694
rect 530506 662660 530910 662692
rect 121458 652176 219562 652286
rect 121458 652112 121532 652176
rect 121596 652112 121632 652176
rect 121696 652112 121734 652176
rect 121798 652112 219562 652176
rect 121458 652080 219562 652112
rect 121458 652016 121530 652080
rect 121594 652016 121632 652080
rect 121696 652016 121730 652080
rect 121794 652016 219562 652080
rect 121458 651886 219562 652016
rect 380992 651018 478142 651116
rect 380992 650954 381064 651018
rect 381128 650954 381164 651018
rect 381228 650954 381266 651018
rect 381330 650954 478142 651018
rect 380992 650922 478142 650954
rect 380992 650858 381062 650922
rect 381126 650858 381164 650922
rect 381228 650858 381262 650922
rect 381326 650858 478142 650922
rect 380992 650716 478142 650858
rect 35278 596592 35923 601996
rect 35277 596454 35924 596592
rect 35277 596218 35506 596454
rect 35742 596218 35924 596454
rect 35277 596134 35924 596218
rect 35277 595898 35506 596134
rect 35742 595928 35924 596134
rect 35742 595898 35925 595928
rect 35277 595856 35925 595898
rect 530510 588794 530910 662660
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 545341 632625 545979 632631
rect 545333 632508 545979 632625
rect 545333 632450 545980 632508
rect 545333 632214 545562 632450
rect 545798 632214 545980 632450
rect 545333 632130 545980 632214
rect 545333 631894 545562 632130
rect 545798 631924 545980 632130
rect 545798 631894 545981 631924
rect 545333 631852 545981 631894
rect 545333 631656 545979 631852
rect 545333 611633 545971 631656
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 545336 597420 545968 611633
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect 545753 578714 546400 585333
rect 545753 578452 546408 578714
rect 545753 578216 545990 578452
rect 546226 578216 546408 578452
rect 545753 578132 546408 578216
rect 545753 577896 545990 578132
rect 546226 577926 546408 578132
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 546226 577896 546409 577926
rect 545753 577854 546409 577896
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 545753 577845 546407 577854
rect 545753 577692 546400 577845
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 530472 475254 530872 475264
rect 530472 475234 530874 475254
rect 530470 475204 530874 475234
rect 530470 475202 530766 475204
rect 530470 475138 530514 475202
rect 530578 475138 530634 475202
rect 530698 475140 530766 475202
rect 530830 475140 530874 475204
rect 530698 475138 530874 475140
rect 530470 475086 530874 475138
rect 530470 475084 530764 475086
rect 530470 475020 530512 475084
rect 530576 475020 530632 475084
rect 530696 475022 530764 475084
rect 530828 475022 530874 475086
rect 530696 475020 530874 475022
rect 530470 474988 530874 475020
rect 530472 474984 530874 474988
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect 34399 470454 35018 470481
rect 34399 470218 34600 470454
rect 34836 470218 35018 470454
rect 34399 470134 35018 470218
rect 34399 469898 34600 470134
rect 34836 469928 35018 470134
rect 34836 469898 35019 469928
rect 34399 469746 35019 469898
rect 34399 442565 35018 469746
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect 34805 416456 35452 430233
rect 34805 416220 35034 416456
rect 35270 416220 35452 416456
rect 34805 416136 35452 416220
rect 34805 415900 35034 416136
rect 35270 415930 35452 416136
rect 35270 415900 35453 415930
rect 34805 415858 35453 415900
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect 49922 351994 50322 436660
rect 530472 404005 530872 474984
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 545331 416446 546006 416568
rect 545331 416210 545560 416446
rect 545796 416210 546006 416446
rect 545331 416126 546006 416210
rect 545331 415890 545560 416126
rect 545796 415890 546006 416126
rect 545331 415740 546006 415890
rect 545339 412437 546006 415740
rect 545722 398652 546373 400601
rect 545720 398518 546373 398652
rect 545720 398460 546374 398518
rect 545720 398224 545956 398460
rect 546192 398224 546374 398460
rect 545720 398140 546374 398224
rect 545720 397904 545956 398140
rect 546192 397934 546374 398140
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 546192 397904 546375 397934
rect 545720 397862 546375 397904
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 545720 397748 546373 397862
rect 49922 351992 50218 351994
rect 49922 351928 49966 351992
rect 50030 351928 50086 351992
rect 50150 351930 50218 351992
rect 50282 351930 50322 351994
rect 50150 351928 50322 351930
rect 49922 351876 50322 351928
rect 49922 351874 50216 351876
rect 49922 351810 49964 351874
rect 50028 351810 50084 351874
rect 50148 351812 50216 351874
rect 50280 351812 50322 351876
rect 50148 351810 50322 351812
rect 49922 351778 50322 351810
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 529338 287568 529738 287592
rect 529336 287548 529738 287568
rect 529332 287518 529738 287548
rect 529332 287516 529628 287518
rect 529332 287452 529376 287516
rect 529440 287452 529496 287516
rect 529560 287454 529628 287516
rect 529692 287454 529738 287518
rect 529560 287452 529738 287454
rect 529332 287400 529738 287452
rect 529332 287398 529626 287400
rect 529332 287334 529374 287398
rect 529438 287334 529494 287398
rect 529558 287336 529626 287398
rect 529690 287336 529738 287400
rect 529558 287334 529738 287336
rect 529332 287302 529738 287334
rect 529336 287292 529738 287302
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect 529338 213778 529738 287292
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 544167 236458 544833 236594
rect 544167 236222 544412 236458
rect 544648 236222 544833 236458
rect 544167 236138 544833 236222
rect 544167 235902 544412 236138
rect 544648 235902 544833 236138
rect 544167 222583 544833 235902
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect 544627 182468 545328 210514
rect 544627 182232 544876 182468
rect 545112 182232 545328 182468
rect 544627 182148 545328 182232
rect 544627 181912 544876 182148
rect 545112 181912 545328 182148
rect 544627 181786 545328 181912
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 18800 -1396 37898
rect -1996 18448 -1814 18800
rect -1506 18448 -1396 18800
rect -1996 17434 -1396 18448
rect -1996 17082 -1812 17434
rect -1504 17082 -1396 17434
rect -1996 15182 -1396 17082
rect -1996 14830 -1850 15182
rect -1542 14830 -1396 15182
rect -1996 2454 -1396 14830
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 -346 1404 480
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 4404 -2226 5004 480
rect 4404 -2462 4586 -2226
rect 4822 -2462 5004 -2226
rect 4404 -2546 5004 -2462
rect 4404 -2782 4586 -2546
rect 4822 -2782 5004 -2546
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 4404 -3744 5004 -2782
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 8004 -4106 8604 480
rect 8004 -4342 8186 -4106
rect 8422 -4342 8604 -4106
rect 8004 -4426 8604 -4342
rect 8004 -4662 8186 -4426
rect 8422 -4662 8604 -4426
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 8004 -5624 8604 -4662
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 11604 -5986 12204 480
rect 18804 -1286 19404 480
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 22404 -3166 23004 480
rect 22404 -3402 22586 -3166
rect 22822 -3402 23004 -3166
rect 22404 -3486 23004 -3402
rect 22404 -3722 22586 -3486
rect 22822 -3722 23004 -3486
rect 22404 -3744 23004 -3722
rect 26004 -5046 26604 480
rect 26004 -5282 26186 -5046
rect 26422 -5282 26604 -5046
rect 26004 -5366 26604 -5282
rect 26004 -5602 26186 -5366
rect 26422 -5602 26604 -5366
rect 26004 -5624 26604 -5602
rect 11604 -6222 11786 -5986
rect 12022 -6222 12204 -5986
rect 11604 -6306 12204 -6222
rect 11604 -6542 11786 -6306
rect 12022 -6542 12204 -6306
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 11604 -7504 12204 -6542
rect 29604 -6926 30204 480
rect 36804 -346 37404 480
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 40404 -2226 41004 480
rect 40404 -2462 40586 -2226
rect 40822 -2462 41004 -2226
rect 40404 -2546 41004 -2462
rect 40404 -2782 40586 -2546
rect 40822 -2782 41004 -2546
rect 40404 -3744 41004 -2782
rect 44004 -4106 44604 480
rect 44004 -4342 44186 -4106
rect 44422 -4342 44604 -4106
rect 44004 -4426 44604 -4342
rect 44004 -4662 44186 -4426
rect 44422 -4662 44604 -4426
rect 44004 -5624 44604 -4662
rect 29604 -7162 29786 -6926
rect 30022 -7162 30204 -6926
rect 29604 -7246 30204 -7162
rect 29604 -7482 29786 -7246
rect 30022 -7482 30204 -7246
rect 29604 -7504 30204 -7482
rect 47604 -5986 48204 480
rect 54804 -1286 55404 480
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 58404 -3166 59004 480
rect 58404 -3402 58586 -3166
rect 58822 -3402 59004 -3166
rect 58404 -3486 59004 -3402
rect 58404 -3722 58586 -3486
rect 58822 -3722 59004 -3486
rect 58404 -3744 59004 -3722
rect 62004 -5046 62604 480
rect 62004 -5282 62186 -5046
rect 62422 -5282 62604 -5046
rect 62004 -5366 62604 -5282
rect 62004 -5602 62186 -5366
rect 62422 -5602 62604 -5366
rect 62004 -5624 62604 -5602
rect 47604 -6222 47786 -5986
rect 48022 -6222 48204 -5986
rect 47604 -6306 48204 -6222
rect 47604 -6542 47786 -6306
rect 48022 -6542 48204 -6306
rect 47604 -7504 48204 -6542
rect 65604 -6926 66204 480
rect 72804 -346 73404 480
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 76404 -2226 77004 480
rect 76404 -2462 76586 -2226
rect 76822 -2462 77004 -2226
rect 76404 -2546 77004 -2462
rect 76404 -2782 76586 -2546
rect 76822 -2782 77004 -2546
rect 76404 -3744 77004 -2782
rect 80004 -4106 80604 480
rect 80004 -4342 80186 -4106
rect 80422 -4342 80604 -4106
rect 80004 -4426 80604 -4342
rect 80004 -4662 80186 -4426
rect 80422 -4662 80604 -4426
rect 80004 -5624 80604 -4662
rect 65604 -7162 65786 -6926
rect 66022 -7162 66204 -6926
rect 65604 -7246 66204 -7162
rect 65604 -7482 65786 -7246
rect 66022 -7482 66204 -7246
rect 65604 -7504 66204 -7482
rect 83604 -5986 84204 480
rect 90804 -1286 91404 480
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 94404 -3166 95004 480
rect 94404 -3402 94586 -3166
rect 94822 -3402 95004 -3166
rect 94404 -3486 95004 -3402
rect 94404 -3722 94586 -3486
rect 94822 -3722 95004 -3486
rect 94404 -3744 95004 -3722
rect 98004 -5046 98604 480
rect 98004 -5282 98186 -5046
rect 98422 -5282 98604 -5046
rect 98004 -5366 98604 -5282
rect 98004 -5602 98186 -5366
rect 98422 -5602 98604 -5366
rect 98004 -5624 98604 -5602
rect 83604 -6222 83786 -5986
rect 84022 -6222 84204 -5986
rect 83604 -6306 84204 -6222
rect 83604 -6542 83786 -6306
rect 84022 -6542 84204 -6306
rect 83604 -7504 84204 -6542
rect 101604 -6926 102204 480
rect 108804 -346 109404 480
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 112404 -2226 113004 480
rect 112404 -2462 112586 -2226
rect 112822 -2462 113004 -2226
rect 112404 -2546 113004 -2462
rect 112404 -2782 112586 -2546
rect 112822 -2782 113004 -2546
rect 112404 -3744 113004 -2782
rect 116004 -4106 116604 480
rect 116004 -4342 116186 -4106
rect 116422 -4342 116604 -4106
rect 116004 -4426 116604 -4342
rect 116004 -4662 116186 -4426
rect 116422 -4662 116604 -4426
rect 116004 -5624 116604 -4662
rect 101604 -7162 101786 -6926
rect 102022 -7162 102204 -6926
rect 101604 -7246 102204 -7162
rect 101604 -7482 101786 -7246
rect 102022 -7482 102204 -7246
rect 101604 -7504 102204 -7482
rect 119604 -5986 120204 480
rect 126804 -1286 127404 480
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 130404 -3166 131004 480
rect 130404 -3402 130586 -3166
rect 130822 -3402 131004 -3166
rect 130404 -3486 131004 -3402
rect 130404 -3722 130586 -3486
rect 130822 -3722 131004 -3486
rect 130404 -3744 131004 -3722
rect 134004 -5046 134604 480
rect 134004 -5282 134186 -5046
rect 134422 -5282 134604 -5046
rect 134004 -5366 134604 -5282
rect 134004 -5602 134186 -5366
rect 134422 -5602 134604 -5366
rect 134004 -5624 134604 -5602
rect 119604 -6222 119786 -5986
rect 120022 -6222 120204 -5986
rect 119604 -6306 120204 -6222
rect 119604 -6542 119786 -6306
rect 120022 -6542 120204 -6306
rect 119604 -7504 120204 -6542
rect 137604 -6926 138204 480
rect 144804 -346 145404 480
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 148404 -2226 149004 480
rect 148404 -2462 148586 -2226
rect 148822 -2462 149004 -2226
rect 148404 -2546 149004 -2462
rect 148404 -2782 148586 -2546
rect 148822 -2782 149004 -2546
rect 148404 -3744 149004 -2782
rect 152004 -4106 152604 480
rect 152004 -4342 152186 -4106
rect 152422 -4342 152604 -4106
rect 152004 -4426 152604 -4342
rect 152004 -4662 152186 -4426
rect 152422 -4662 152604 -4426
rect 152004 -5624 152604 -4662
rect 137604 -7162 137786 -6926
rect 138022 -7162 138204 -6926
rect 137604 -7246 138204 -7162
rect 137604 -7482 137786 -7246
rect 138022 -7482 138204 -7246
rect 137604 -7504 138204 -7482
rect 155604 -5986 156204 480
rect 162804 -1286 163404 480
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 166404 -3166 167004 480
rect 166404 -3402 166586 -3166
rect 166822 -3402 167004 -3166
rect 166404 -3486 167004 -3402
rect 166404 -3722 166586 -3486
rect 166822 -3722 167004 -3486
rect 166404 -3744 167004 -3722
rect 170004 -5046 170604 480
rect 170004 -5282 170186 -5046
rect 170422 -5282 170604 -5046
rect 170004 -5366 170604 -5282
rect 170004 -5602 170186 -5366
rect 170422 -5602 170604 -5366
rect 170004 -5624 170604 -5602
rect 155604 -6222 155786 -5986
rect 156022 -6222 156204 -5986
rect 155604 -6306 156204 -6222
rect 155604 -6542 155786 -6306
rect 156022 -6542 156204 -6306
rect 155604 -7504 156204 -6542
rect 173604 -6926 174204 480
rect 180804 -346 181404 480
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 184404 -2226 185004 480
rect 184404 -2462 184586 -2226
rect 184822 -2462 185004 -2226
rect 184404 -2546 185004 -2462
rect 184404 -2782 184586 -2546
rect 184822 -2782 185004 -2546
rect 184404 -3744 185004 -2782
rect 188004 -4106 188604 480
rect 188004 -4342 188186 -4106
rect 188422 -4342 188604 -4106
rect 188004 -4426 188604 -4342
rect 188004 -4662 188186 -4426
rect 188422 -4662 188604 -4426
rect 188004 -5624 188604 -4662
rect 173604 -7162 173786 -6926
rect 174022 -7162 174204 -6926
rect 173604 -7246 174204 -7162
rect 173604 -7482 173786 -7246
rect 174022 -7482 174204 -7246
rect 173604 -7504 174204 -7482
rect 191604 -5986 192204 480
rect 198804 -1286 199404 480
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 202404 -3166 203004 480
rect 202404 -3402 202586 -3166
rect 202822 -3402 203004 -3166
rect 202404 -3486 203004 -3402
rect 202404 -3722 202586 -3486
rect 202822 -3722 203004 -3486
rect 202404 -3744 203004 -3722
rect 206004 -5046 206604 480
rect 206004 -5282 206186 -5046
rect 206422 -5282 206604 -5046
rect 206004 -5366 206604 -5282
rect 206004 -5602 206186 -5366
rect 206422 -5602 206604 -5366
rect 206004 -5624 206604 -5602
rect 191604 -6222 191786 -5986
rect 192022 -6222 192204 -5986
rect 191604 -6306 192204 -6222
rect 191604 -6542 191786 -6306
rect 192022 -6542 192204 -6306
rect 191604 -7504 192204 -6542
rect 209604 -6926 210204 480
rect 216804 -346 217404 480
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 220404 -2226 221004 480
rect 220404 -2462 220586 -2226
rect 220822 -2462 221004 -2226
rect 220404 -2546 221004 -2462
rect 220404 -2782 220586 -2546
rect 220822 -2782 221004 -2546
rect 220404 -3744 221004 -2782
rect 224004 -4106 224604 480
rect 224004 -4342 224186 -4106
rect 224422 -4342 224604 -4106
rect 224004 -4426 224604 -4342
rect 224004 -4662 224186 -4426
rect 224422 -4662 224604 -4426
rect 224004 -5624 224604 -4662
rect 209604 -7162 209786 -6926
rect 210022 -7162 210204 -6926
rect 209604 -7246 210204 -7162
rect 209604 -7482 209786 -7246
rect 210022 -7482 210204 -7246
rect 209604 -7504 210204 -7482
rect 227604 -5986 228204 480
rect 234804 -1286 235404 480
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 238404 -3166 239004 480
rect 238404 -3402 238586 -3166
rect 238822 -3402 239004 -3166
rect 238404 -3486 239004 -3402
rect 238404 -3722 238586 -3486
rect 238822 -3722 239004 -3486
rect 238404 -3744 239004 -3722
rect 242004 -5046 242604 480
rect 242004 -5282 242186 -5046
rect 242422 -5282 242604 -5046
rect 242004 -5366 242604 -5282
rect 242004 -5602 242186 -5366
rect 242422 -5602 242604 -5366
rect 242004 -5624 242604 -5602
rect 227604 -6222 227786 -5986
rect 228022 -6222 228204 -5986
rect 227604 -6306 228204 -6222
rect 227604 -6542 227786 -6306
rect 228022 -6542 228204 -6306
rect 227604 -7504 228204 -6542
rect 245604 -6926 246204 480
rect 252804 -346 253404 480
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 256404 -2226 257004 480
rect 256404 -2462 256586 -2226
rect 256822 -2462 257004 -2226
rect 256404 -2546 257004 -2462
rect 256404 -2782 256586 -2546
rect 256822 -2782 257004 -2546
rect 256404 -3744 257004 -2782
rect 260004 -4106 260604 480
rect 260004 -4342 260186 -4106
rect 260422 -4342 260604 -4106
rect 260004 -4426 260604 -4342
rect 260004 -4662 260186 -4426
rect 260422 -4662 260604 -4426
rect 260004 -5624 260604 -4662
rect 245604 -7162 245786 -6926
rect 246022 -7162 246204 -6926
rect 245604 -7246 246204 -7162
rect 245604 -7482 245786 -7246
rect 246022 -7482 246204 -7246
rect 245604 -7504 246204 -7482
rect 263604 -5986 264204 480
rect 270804 -1286 271404 480
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 274404 -3166 275004 480
rect 274404 -3402 274586 -3166
rect 274822 -3402 275004 -3166
rect 274404 -3486 275004 -3402
rect 274404 -3722 274586 -3486
rect 274822 -3722 275004 -3486
rect 274404 -3744 275004 -3722
rect 278004 -5046 278604 480
rect 278004 -5282 278186 -5046
rect 278422 -5282 278604 -5046
rect 278004 -5366 278604 -5282
rect 278004 -5602 278186 -5366
rect 278422 -5602 278604 -5366
rect 278004 -5624 278604 -5602
rect 263604 -6222 263786 -5986
rect 264022 -6222 264204 -5986
rect 263604 -6306 264204 -6222
rect 263604 -6542 263786 -6306
rect 264022 -6542 264204 -6306
rect 263604 -7504 264204 -6542
rect 281604 -6926 282204 480
rect 288804 -346 289404 480
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 292404 -2226 293004 480
rect 292404 -2462 292586 -2226
rect 292822 -2462 293004 -2226
rect 292404 -2546 293004 -2462
rect 292404 -2782 292586 -2546
rect 292822 -2782 293004 -2546
rect 292404 -3744 293004 -2782
rect 296004 -4106 296604 480
rect 296004 -4342 296186 -4106
rect 296422 -4342 296604 -4106
rect 296004 -4426 296604 -4342
rect 296004 -4662 296186 -4426
rect 296422 -4662 296604 -4426
rect 296004 -5624 296604 -4662
rect 281604 -7162 281786 -6926
rect 282022 -7162 282204 -6926
rect 281604 -7246 282204 -7162
rect 281604 -7482 281786 -7246
rect 282022 -7482 282204 -7246
rect 281604 -7504 282204 -7482
rect 299604 -5986 300204 480
rect 306804 -1286 307404 480
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 310404 -3166 311004 480
rect 310404 -3402 310586 -3166
rect 310822 -3402 311004 -3166
rect 310404 -3486 311004 -3402
rect 310404 -3722 310586 -3486
rect 310822 -3722 311004 -3486
rect 310404 -3744 311004 -3722
rect 314004 -5046 314604 480
rect 314004 -5282 314186 -5046
rect 314422 -5282 314604 -5046
rect 314004 -5366 314604 -5282
rect 314004 -5602 314186 -5366
rect 314422 -5602 314604 -5366
rect 314004 -5624 314604 -5602
rect 299604 -6222 299786 -5986
rect 300022 -6222 300204 -5986
rect 299604 -6306 300204 -6222
rect 299604 -6542 299786 -6306
rect 300022 -6542 300204 -6306
rect 299604 -7504 300204 -6542
rect 317604 -6926 318204 480
rect 324804 -346 325404 480
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 328404 -2226 329004 480
rect 328404 -2462 328586 -2226
rect 328822 -2462 329004 -2226
rect 328404 -2546 329004 -2462
rect 328404 -2782 328586 -2546
rect 328822 -2782 329004 -2546
rect 328404 -3744 329004 -2782
rect 332004 -4106 332604 480
rect 332004 -4342 332186 -4106
rect 332422 -4342 332604 -4106
rect 332004 -4426 332604 -4342
rect 332004 -4662 332186 -4426
rect 332422 -4662 332604 -4426
rect 332004 -5624 332604 -4662
rect 317604 -7162 317786 -6926
rect 318022 -7162 318204 -6926
rect 317604 -7246 318204 -7162
rect 317604 -7482 317786 -7246
rect 318022 -7482 318204 -7246
rect 317604 -7504 318204 -7482
rect 335604 -5986 336204 480
rect 342804 -1286 343404 480
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 346404 -3166 347004 480
rect 346404 -3402 346586 -3166
rect 346822 -3402 347004 -3166
rect 346404 -3486 347004 -3402
rect 346404 -3722 346586 -3486
rect 346822 -3722 347004 -3486
rect 346404 -3744 347004 -3722
rect 350004 -5046 350604 480
rect 350004 -5282 350186 -5046
rect 350422 -5282 350604 -5046
rect 350004 -5366 350604 -5282
rect 350004 -5602 350186 -5366
rect 350422 -5602 350604 -5366
rect 350004 -5624 350604 -5602
rect 335604 -6222 335786 -5986
rect 336022 -6222 336204 -5986
rect 335604 -6306 336204 -6222
rect 335604 -6542 335786 -6306
rect 336022 -6542 336204 -6306
rect 335604 -7504 336204 -6542
rect 353604 -6926 354204 480
rect 360804 -346 361404 480
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 364404 -2226 365004 480
rect 364404 -2462 364586 -2226
rect 364822 -2462 365004 -2226
rect 364404 -2546 365004 -2462
rect 364404 -2782 364586 -2546
rect 364822 -2782 365004 -2546
rect 364404 -3744 365004 -2782
rect 368004 -4106 368604 480
rect 368004 -4342 368186 -4106
rect 368422 -4342 368604 -4106
rect 368004 -4426 368604 -4342
rect 368004 -4662 368186 -4426
rect 368422 -4662 368604 -4426
rect 368004 -5624 368604 -4662
rect 353604 -7162 353786 -6926
rect 354022 -7162 354204 -6926
rect 353604 -7246 354204 -7162
rect 353604 -7482 353786 -7246
rect 354022 -7482 354204 -7246
rect 353604 -7504 354204 -7482
rect 371604 -5986 372204 480
rect 378804 -1286 379404 480
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 382404 -3166 383004 480
rect 382404 -3402 382586 -3166
rect 382822 -3402 383004 -3166
rect 382404 -3486 383004 -3402
rect 382404 -3722 382586 -3486
rect 382822 -3722 383004 -3486
rect 382404 -3744 383004 -3722
rect 386004 -5046 386604 480
rect 386004 -5282 386186 -5046
rect 386422 -5282 386604 -5046
rect 386004 -5366 386604 -5282
rect 386004 -5602 386186 -5366
rect 386422 -5602 386604 -5366
rect 386004 -5624 386604 -5602
rect 371604 -6222 371786 -5986
rect 372022 -6222 372204 -5986
rect 371604 -6306 372204 -6222
rect 371604 -6542 371786 -6306
rect 372022 -6542 372204 -6306
rect 371604 -7504 372204 -6542
rect 389604 -6926 390204 480
rect 396804 -346 397404 480
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 400404 -2226 401004 480
rect 400404 -2462 400586 -2226
rect 400822 -2462 401004 -2226
rect 400404 -2546 401004 -2462
rect 400404 -2782 400586 -2546
rect 400822 -2782 401004 -2546
rect 400404 -3744 401004 -2782
rect 404004 -4106 404604 480
rect 404004 -4342 404186 -4106
rect 404422 -4342 404604 -4106
rect 404004 -4426 404604 -4342
rect 404004 -4662 404186 -4426
rect 404422 -4662 404604 -4426
rect 404004 -5624 404604 -4662
rect 389604 -7162 389786 -6926
rect 390022 -7162 390204 -6926
rect 389604 -7246 390204 -7162
rect 389604 -7482 389786 -7246
rect 390022 -7482 390204 -7246
rect 389604 -7504 390204 -7482
rect 407604 -5986 408204 480
rect 414804 -1286 415404 480
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 418404 -3166 419004 480
rect 418404 -3402 418586 -3166
rect 418822 -3402 419004 -3166
rect 418404 -3486 419004 -3402
rect 418404 -3722 418586 -3486
rect 418822 -3722 419004 -3486
rect 418404 -3744 419004 -3722
rect 422004 -5046 422604 480
rect 422004 -5282 422186 -5046
rect 422422 -5282 422604 -5046
rect 422004 -5366 422604 -5282
rect 422004 -5602 422186 -5366
rect 422422 -5602 422604 -5366
rect 422004 -5624 422604 -5602
rect 407604 -6222 407786 -5986
rect 408022 -6222 408204 -5986
rect 407604 -6306 408204 -6222
rect 407604 -6542 407786 -6306
rect 408022 -6542 408204 -6306
rect 407604 -7504 408204 -6542
rect 425604 -6926 426204 480
rect 432804 -346 433404 480
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 436404 -2226 437004 480
rect 436404 -2462 436586 -2226
rect 436822 -2462 437004 -2226
rect 436404 -2546 437004 -2462
rect 436404 -2782 436586 -2546
rect 436822 -2782 437004 -2546
rect 436404 -3744 437004 -2782
rect 440004 -4106 440604 480
rect 440004 -4342 440186 -4106
rect 440422 -4342 440604 -4106
rect 440004 -4426 440604 -4342
rect 440004 -4662 440186 -4426
rect 440422 -4662 440604 -4426
rect 440004 -5624 440604 -4662
rect 425604 -7162 425786 -6926
rect 426022 -7162 426204 -6926
rect 425604 -7246 426204 -7162
rect 425604 -7482 425786 -7246
rect 426022 -7482 426204 -7246
rect 425604 -7504 426204 -7482
rect 443604 -5986 444204 480
rect 450804 -1286 451404 480
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 454404 -3166 455004 480
rect 454404 -3402 454586 -3166
rect 454822 -3402 455004 -3166
rect 454404 -3486 455004 -3402
rect 454404 -3722 454586 -3486
rect 454822 -3722 455004 -3486
rect 454404 -3744 455004 -3722
rect 458004 -5046 458604 480
rect 458004 -5282 458186 -5046
rect 458422 -5282 458604 -5046
rect 458004 -5366 458604 -5282
rect 458004 -5602 458186 -5366
rect 458422 -5602 458604 -5366
rect 458004 -5624 458604 -5602
rect 443604 -6222 443786 -5986
rect 444022 -6222 444204 -5986
rect 443604 -6306 444204 -6222
rect 443604 -6542 443786 -6306
rect 444022 -6542 444204 -6306
rect 443604 -7504 444204 -6542
rect 461604 -6926 462204 480
rect 468804 -346 469404 480
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 472404 -2226 473004 480
rect 472404 -2462 472586 -2226
rect 472822 -2462 473004 -2226
rect 472404 -2546 473004 -2462
rect 472404 -2782 472586 -2546
rect 472822 -2782 473004 -2546
rect 472404 -3744 473004 -2782
rect 476004 -4106 476604 480
rect 476004 -4342 476186 -4106
rect 476422 -4342 476604 -4106
rect 476004 -4426 476604 -4342
rect 476004 -4662 476186 -4426
rect 476422 -4662 476604 -4426
rect 476004 -5624 476604 -4662
rect 461604 -7162 461786 -6926
rect 462022 -7162 462204 -6926
rect 461604 -7246 462204 -7162
rect 461604 -7482 461786 -7246
rect 462022 -7482 462204 -7246
rect 461604 -7504 462204 -7482
rect 479604 -5986 480204 480
rect 486804 -1286 487404 480
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 490404 -3166 491004 480
rect 490404 -3402 490586 -3166
rect 490822 -3402 491004 -3166
rect 490404 -3486 491004 -3402
rect 490404 -3722 490586 -3486
rect 490822 -3722 491004 -3486
rect 490404 -3744 491004 -3722
rect 494004 -5046 494604 480
rect 494004 -5282 494186 -5046
rect 494422 -5282 494604 -5046
rect 494004 -5366 494604 -5282
rect 494004 -5602 494186 -5366
rect 494422 -5602 494604 -5366
rect 494004 -5624 494604 -5602
rect 479604 -6222 479786 -5986
rect 480022 -6222 480204 -5986
rect 479604 -6306 480204 -6222
rect 479604 -6542 479786 -6306
rect 480022 -6542 480204 -6306
rect 479604 -7504 480204 -6542
rect 497604 -6926 498204 480
rect 504804 -346 505404 480
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 508404 -2226 509004 480
rect 508404 -2462 508586 -2226
rect 508822 -2462 509004 -2226
rect 508404 -2546 509004 -2462
rect 508404 -2782 508586 -2546
rect 508822 -2782 509004 -2546
rect 508404 -3744 509004 -2782
rect 512004 -4106 512604 480
rect 512004 -4342 512186 -4106
rect 512422 -4342 512604 -4106
rect 512004 -4426 512604 -4342
rect 512004 -4662 512186 -4426
rect 512422 -4662 512604 -4426
rect 512004 -5624 512604 -4662
rect 497604 -7162 497786 -6926
rect 498022 -7162 498204 -6926
rect 497604 -7246 498204 -7162
rect 497604 -7482 497786 -7246
rect 498022 -7482 498204 -7246
rect 497604 -7504 498204 -7482
rect 515604 -5986 516204 480
rect 522804 -1286 523404 480
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 526404 -3166 527004 480
rect 526404 -3402 526586 -3166
rect 526822 -3402 527004 -3166
rect 526404 -3486 527004 -3402
rect 526404 -3722 526586 -3486
rect 526822 -3722 527004 -3486
rect 526404 -3744 527004 -3722
rect 530004 -5046 530604 480
rect 530004 -5282 530186 -5046
rect 530422 -5282 530604 -5046
rect 530004 -5366 530604 -5282
rect 530004 -5602 530186 -5366
rect 530422 -5602 530604 -5366
rect 530004 -5624 530604 -5602
rect 515604 -6222 515786 -5986
rect 516022 -6222 516204 -5986
rect 515604 -6306 516204 -6222
rect 515604 -6542 515786 -6306
rect 516022 -6542 516204 -6306
rect 515604 -7504 516204 -6542
rect 533604 -6926 534204 480
rect 540804 -346 541404 480
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 544404 -2226 545004 480
rect 544404 -2462 544586 -2226
rect 544822 -2462 545004 -2226
rect 544404 -2546 545004 -2462
rect 544404 -2782 544586 -2546
rect 544822 -2782 545004 -2546
rect 544404 -3744 545004 -2782
rect 548004 -4106 548604 480
rect 548004 -4342 548186 -4106
rect 548422 -4342 548604 -4106
rect 548004 -4426 548604 -4342
rect 548004 -4662 548186 -4426
rect 548422 -4662 548604 -4426
rect 548004 -5624 548604 -4662
rect 533604 -7162 533786 -6926
rect 534022 -7162 534204 -6926
rect 533604 -7246 534204 -7162
rect 533604 -7482 533786 -7246
rect 534022 -7482 534204 -7246
rect 533604 -7504 534204 -7482
rect 551604 -5986 552204 480
rect 558804 -1286 559404 480
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 562404 -3166 563004 480
rect 562404 -3402 562586 -3166
rect 562822 -3402 563004 -3166
rect 562404 -3486 563004 -3402
rect 562404 -3722 562586 -3486
rect 562822 -3722 563004 -3486
rect 562404 -3744 563004 -3722
rect 566004 -5046 566604 480
rect 566004 -5282 566186 -5046
rect 566422 -5282 566604 -5046
rect 566004 -5366 566604 -5282
rect 566004 -5602 566186 -5366
rect 566422 -5602 566604 -5366
rect 566004 -5624 566604 -5602
rect 551604 -6222 551786 -5986
rect 552022 -6222 552204 -5986
rect 551604 -6306 552204 -6222
rect 551604 -6542 551786 -6306
rect 552022 -6542 552204 -6306
rect 551604 -7504 552204 -6542
rect 569604 -6926 570204 480
rect 576804 -346 577404 480
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 580404 -2226 581004 480
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 587200 690054 587800 706162
rect 587200 689818 587382 690054
rect 587618 689818 587800 690054
rect 587200 689734 587800 689818
rect 587200 689498 587382 689734
rect 587618 689498 587800 689734
rect 587200 654054 587800 689498
rect 587200 653818 587382 654054
rect 587618 653818 587800 654054
rect 587200 653734 587800 653818
rect 587200 653498 587382 653734
rect 587618 653498 587800 653734
rect 587200 618054 587800 653498
rect 587200 617818 587382 618054
rect 587618 617818 587800 618054
rect 587200 617734 587800 617818
rect 587200 617498 587382 617734
rect 587618 617498 587800 617734
rect 587200 582054 587800 617498
rect 587200 581818 587382 582054
rect 587618 581818 587800 582054
rect 587200 581734 587800 581818
rect 587200 581498 587382 581734
rect 587618 581498 587800 581734
rect 587200 546054 587800 581498
rect 587200 545818 587382 546054
rect 587618 545818 587800 546054
rect 587200 545734 587800 545818
rect 587200 545498 587382 545734
rect 587618 545498 587800 545734
rect 587200 510054 587800 545498
rect 587200 509818 587382 510054
rect 587618 509818 587800 510054
rect 587200 509734 587800 509818
rect 587200 509498 587382 509734
rect 587618 509498 587800 509734
rect 587200 474054 587800 509498
rect 587200 473818 587382 474054
rect 587618 473818 587800 474054
rect 587200 473734 587800 473818
rect 587200 473498 587382 473734
rect 587618 473498 587800 473734
rect 587200 438054 587800 473498
rect 587200 437818 587382 438054
rect 587618 437818 587800 438054
rect 587200 437734 587800 437818
rect 587200 437498 587382 437734
rect 587618 437498 587800 437734
rect 587200 402054 587800 437498
rect 587200 401818 587382 402054
rect 587618 401818 587800 402054
rect 587200 401734 587800 401818
rect 587200 401498 587382 401734
rect 587618 401498 587800 401734
rect 587200 366054 587800 401498
rect 587200 365818 587382 366054
rect 587618 365818 587800 366054
rect 587200 365734 587800 365818
rect 587200 365498 587382 365734
rect 587618 365498 587800 365734
rect 587200 330054 587800 365498
rect 587200 329818 587382 330054
rect 587618 329818 587800 330054
rect 587200 329734 587800 329818
rect 587200 329498 587382 329734
rect 587618 329498 587800 329734
rect 587200 294054 587800 329498
rect 587200 293818 587382 294054
rect 587618 293818 587800 294054
rect 587200 293734 587800 293818
rect 587200 293498 587382 293734
rect 587618 293498 587800 293734
rect 587200 258054 587800 293498
rect 587200 257818 587382 258054
rect 587618 257818 587800 258054
rect 587200 257734 587800 257818
rect 587200 257498 587382 257734
rect 587618 257498 587800 257734
rect 587200 222054 587800 257498
rect 587200 221818 587382 222054
rect 587618 221818 587800 222054
rect 587200 221734 587800 221818
rect 587200 221498 587382 221734
rect 587618 221498 587800 221734
rect 587200 186054 587800 221498
rect 587200 185818 587382 186054
rect 587618 185818 587800 186054
rect 587200 185734 587800 185818
rect 587200 185498 587382 185734
rect 587618 185498 587800 185734
rect 587200 150054 587800 185498
rect 587200 149818 587382 150054
rect 587618 149818 587800 150054
rect 587200 149734 587800 149818
rect 587200 149498 587382 149734
rect 587618 149498 587800 149734
rect 587200 114054 587800 149498
rect 587200 113818 587382 114054
rect 587618 113818 587800 114054
rect 587200 113734 587800 113818
rect 587200 113498 587382 113734
rect 587618 113498 587800 113734
rect 587200 78054 587800 113498
rect 587200 77818 587382 78054
rect 587618 77818 587800 78054
rect 587200 77734 587800 77818
rect 587200 77498 587382 77734
rect 587618 77498 587800 77734
rect 587200 42054 587800 77498
rect 587200 41818 587382 42054
rect 587618 41818 587800 42054
rect 587200 41734 587800 41818
rect 587200 41498 587382 41734
rect 587618 41498 587800 41734
rect 587200 6054 587800 41498
rect 587200 5818 587382 6054
rect 587618 5818 587800 6054
rect 587200 5734 587800 5818
rect 587200 5498 587382 5734
rect 587618 5498 587800 5734
rect 580404 -2462 580586 -2226
rect 580822 -2462 581004 -2226
rect 580404 -2546 581004 -2462
rect 580404 -2782 580586 -2546
rect 580822 -2782 581004 -2546
rect 580404 -3744 581004 -2782
rect 587200 -2226 587800 5498
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 672054 588740 707102
rect 588140 671818 588322 672054
rect 588558 671818 588740 672054
rect 588140 671734 588740 671818
rect 588140 671498 588322 671734
rect 588558 671498 588740 671734
rect 588140 636054 588740 671498
rect 588140 635818 588322 636054
rect 588558 635818 588740 636054
rect 588140 635734 588740 635818
rect 588140 635498 588322 635734
rect 588558 635498 588740 635734
rect 588140 600054 588740 635498
rect 588140 599818 588322 600054
rect 588558 599818 588740 600054
rect 588140 599734 588740 599818
rect 588140 599498 588322 599734
rect 588558 599498 588740 599734
rect 588140 564054 588740 599498
rect 588140 563818 588322 564054
rect 588558 563818 588740 564054
rect 588140 563734 588740 563818
rect 588140 563498 588322 563734
rect 588558 563498 588740 563734
rect 588140 528054 588740 563498
rect 588140 527818 588322 528054
rect 588558 527818 588740 528054
rect 588140 527734 588740 527818
rect 588140 527498 588322 527734
rect 588558 527498 588740 527734
rect 588140 492054 588740 527498
rect 588140 491818 588322 492054
rect 588558 491818 588740 492054
rect 588140 491734 588740 491818
rect 588140 491498 588322 491734
rect 588558 491498 588740 491734
rect 588140 456054 588740 491498
rect 588140 455818 588322 456054
rect 588558 455818 588740 456054
rect 588140 455734 588740 455818
rect 588140 455498 588322 455734
rect 588558 455498 588740 455734
rect 588140 420054 588740 455498
rect 588140 419818 588322 420054
rect 588558 419818 588740 420054
rect 588140 419734 588740 419818
rect 588140 419498 588322 419734
rect 588558 419498 588740 419734
rect 588140 384054 588740 419498
rect 588140 383818 588322 384054
rect 588558 383818 588740 384054
rect 588140 383734 588740 383818
rect 588140 383498 588322 383734
rect 588558 383498 588740 383734
rect 588140 348054 588740 383498
rect 588140 347818 588322 348054
rect 588558 347818 588740 348054
rect 588140 347734 588740 347818
rect 588140 347498 588322 347734
rect 588558 347498 588740 347734
rect 588140 312054 588740 347498
rect 588140 311818 588322 312054
rect 588558 311818 588740 312054
rect 588140 311734 588740 311818
rect 588140 311498 588322 311734
rect 588558 311498 588740 311734
rect 588140 276054 588740 311498
rect 588140 275818 588322 276054
rect 588558 275818 588740 276054
rect 588140 275734 588740 275818
rect 588140 275498 588322 275734
rect 588558 275498 588740 275734
rect 588140 240054 588740 275498
rect 588140 239818 588322 240054
rect 588558 239818 588740 240054
rect 588140 239734 588740 239818
rect 588140 239498 588322 239734
rect 588558 239498 588740 239734
rect 588140 204054 588740 239498
rect 588140 203818 588322 204054
rect 588558 203818 588740 204054
rect 588140 203734 588740 203818
rect 588140 203498 588322 203734
rect 588558 203498 588740 203734
rect 588140 168054 588740 203498
rect 588140 167818 588322 168054
rect 588558 167818 588740 168054
rect 588140 167734 588740 167818
rect 588140 167498 588322 167734
rect 588558 167498 588740 167734
rect 588140 132054 588740 167498
rect 588140 131818 588322 132054
rect 588558 131818 588740 132054
rect 588140 131734 588740 131818
rect 588140 131498 588322 131734
rect 588558 131498 588740 131734
rect 588140 96054 588740 131498
rect 588140 95818 588322 96054
rect 588558 95818 588740 96054
rect 588140 95734 588740 95818
rect 588140 95498 588322 95734
rect 588558 95498 588740 95734
rect 588140 60054 588740 95498
rect 588140 59818 588322 60054
rect 588558 59818 588740 60054
rect 588140 59734 588740 59818
rect 588140 59498 588322 59734
rect 588558 59498 588740 59734
rect 588140 24054 588740 59498
rect 588140 23818 588322 24054
rect 588558 23818 588740 24054
rect 588140 23734 588740 23818
rect 588140 23498 588322 23734
rect 588558 23498 588740 23734
rect 588140 -3166 588740 23498
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect 589080 693654 589680 708042
rect 589080 693418 589262 693654
rect 589498 693418 589680 693654
rect 589080 693334 589680 693418
rect 589080 693098 589262 693334
rect 589498 693098 589680 693334
rect 589080 657654 589680 693098
rect 589080 657418 589262 657654
rect 589498 657418 589680 657654
rect 589080 657334 589680 657418
rect 589080 657098 589262 657334
rect 589498 657098 589680 657334
rect 589080 621654 589680 657098
rect 589080 621418 589262 621654
rect 589498 621418 589680 621654
rect 589080 621334 589680 621418
rect 589080 621098 589262 621334
rect 589498 621098 589680 621334
rect 589080 585654 589680 621098
rect 589080 585418 589262 585654
rect 589498 585418 589680 585654
rect 589080 585334 589680 585418
rect 589080 585098 589262 585334
rect 589498 585098 589680 585334
rect 589080 549654 589680 585098
rect 589080 549418 589262 549654
rect 589498 549418 589680 549654
rect 589080 549334 589680 549418
rect 589080 549098 589262 549334
rect 589498 549098 589680 549334
rect 589080 513654 589680 549098
rect 589080 513418 589262 513654
rect 589498 513418 589680 513654
rect 589080 513334 589680 513418
rect 589080 513098 589262 513334
rect 589498 513098 589680 513334
rect 589080 477654 589680 513098
rect 589080 477418 589262 477654
rect 589498 477418 589680 477654
rect 589080 477334 589680 477418
rect 589080 477098 589262 477334
rect 589498 477098 589680 477334
rect 589080 441654 589680 477098
rect 589080 441418 589262 441654
rect 589498 441418 589680 441654
rect 589080 441334 589680 441418
rect 589080 441098 589262 441334
rect 589498 441098 589680 441334
rect 589080 405654 589680 441098
rect 589080 405418 589262 405654
rect 589498 405418 589680 405654
rect 589080 405334 589680 405418
rect 589080 405098 589262 405334
rect 589498 405098 589680 405334
rect 589080 369654 589680 405098
rect 589080 369418 589262 369654
rect 589498 369418 589680 369654
rect 589080 369334 589680 369418
rect 589080 369098 589262 369334
rect 589498 369098 589680 369334
rect 589080 333654 589680 369098
rect 589080 333418 589262 333654
rect 589498 333418 589680 333654
rect 589080 333334 589680 333418
rect 589080 333098 589262 333334
rect 589498 333098 589680 333334
rect 589080 297654 589680 333098
rect 589080 297418 589262 297654
rect 589498 297418 589680 297654
rect 589080 297334 589680 297418
rect 589080 297098 589262 297334
rect 589498 297098 589680 297334
rect 589080 261654 589680 297098
rect 589080 261418 589262 261654
rect 589498 261418 589680 261654
rect 589080 261334 589680 261418
rect 589080 261098 589262 261334
rect 589498 261098 589680 261334
rect 589080 225654 589680 261098
rect 589080 225418 589262 225654
rect 589498 225418 589680 225654
rect 589080 225334 589680 225418
rect 589080 225098 589262 225334
rect 589498 225098 589680 225334
rect 589080 189654 589680 225098
rect 589080 189418 589262 189654
rect 589498 189418 589680 189654
rect 589080 189334 589680 189418
rect 589080 189098 589262 189334
rect 589498 189098 589680 189334
rect 589080 153654 589680 189098
rect 589080 153418 589262 153654
rect 589498 153418 589680 153654
rect 589080 153334 589680 153418
rect 589080 153098 589262 153334
rect 589498 153098 589680 153334
rect 589080 117654 589680 153098
rect 589080 117418 589262 117654
rect 589498 117418 589680 117654
rect 589080 117334 589680 117418
rect 589080 117098 589262 117334
rect 589498 117098 589680 117334
rect 589080 81654 589680 117098
rect 589080 81418 589262 81654
rect 589498 81418 589680 81654
rect 589080 81334 589680 81418
rect 589080 81098 589262 81334
rect 589498 81098 589680 81334
rect 589080 45654 589680 81098
rect 589080 45418 589262 45654
rect 589498 45418 589680 45654
rect 589080 45334 589680 45418
rect 589080 45098 589262 45334
rect 589498 45098 589680 45334
rect 589080 9654 589680 45098
rect 589080 9418 589262 9654
rect 589498 9418 589680 9654
rect 589080 9334 589680 9418
rect 589080 9098 589262 9334
rect 589498 9098 589680 9334
rect 589080 -4106 589680 9098
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect 590020 675654 590620 708982
rect 590020 675418 590202 675654
rect 590438 675418 590620 675654
rect 590020 675334 590620 675418
rect 590020 675098 590202 675334
rect 590438 675098 590620 675334
rect 590020 639654 590620 675098
rect 590020 639418 590202 639654
rect 590438 639418 590620 639654
rect 590020 639334 590620 639418
rect 590020 639098 590202 639334
rect 590438 639098 590620 639334
rect 590020 603654 590620 639098
rect 590020 603418 590202 603654
rect 590438 603418 590620 603654
rect 590020 603334 590620 603418
rect 590020 603098 590202 603334
rect 590438 603098 590620 603334
rect 590020 567654 590620 603098
rect 590020 567418 590202 567654
rect 590438 567418 590620 567654
rect 590020 567334 590620 567418
rect 590020 567098 590202 567334
rect 590438 567098 590620 567334
rect 590020 531654 590620 567098
rect 590020 531418 590202 531654
rect 590438 531418 590620 531654
rect 590020 531334 590620 531418
rect 590020 531098 590202 531334
rect 590438 531098 590620 531334
rect 590020 495654 590620 531098
rect 590020 495418 590202 495654
rect 590438 495418 590620 495654
rect 590020 495334 590620 495418
rect 590020 495098 590202 495334
rect 590438 495098 590620 495334
rect 590020 459654 590620 495098
rect 590020 459418 590202 459654
rect 590438 459418 590620 459654
rect 590020 459334 590620 459418
rect 590020 459098 590202 459334
rect 590438 459098 590620 459334
rect 590020 423654 590620 459098
rect 590020 423418 590202 423654
rect 590438 423418 590620 423654
rect 590020 423334 590620 423418
rect 590020 423098 590202 423334
rect 590438 423098 590620 423334
rect 590020 387654 590620 423098
rect 590020 387418 590202 387654
rect 590438 387418 590620 387654
rect 590020 387334 590620 387418
rect 590020 387098 590202 387334
rect 590438 387098 590620 387334
rect 590020 351654 590620 387098
rect 590020 351418 590202 351654
rect 590438 351418 590620 351654
rect 590020 351334 590620 351418
rect 590020 351098 590202 351334
rect 590438 351098 590620 351334
rect 590020 315654 590620 351098
rect 590020 315418 590202 315654
rect 590438 315418 590620 315654
rect 590020 315334 590620 315418
rect 590020 315098 590202 315334
rect 590438 315098 590620 315334
rect 590020 279654 590620 315098
rect 590020 279418 590202 279654
rect 590438 279418 590620 279654
rect 590020 279334 590620 279418
rect 590020 279098 590202 279334
rect 590438 279098 590620 279334
rect 590020 243654 590620 279098
rect 590020 243418 590202 243654
rect 590438 243418 590620 243654
rect 590020 243334 590620 243418
rect 590020 243098 590202 243334
rect 590438 243098 590620 243334
rect 590020 207654 590620 243098
rect 590020 207418 590202 207654
rect 590438 207418 590620 207654
rect 590020 207334 590620 207418
rect 590020 207098 590202 207334
rect 590438 207098 590620 207334
rect 590020 171654 590620 207098
rect 590020 171418 590202 171654
rect 590438 171418 590620 171654
rect 590020 171334 590620 171418
rect 590020 171098 590202 171334
rect 590438 171098 590620 171334
rect 590020 135654 590620 171098
rect 590020 135418 590202 135654
rect 590438 135418 590620 135654
rect 590020 135334 590620 135418
rect 590020 135098 590202 135334
rect 590438 135098 590620 135334
rect 590020 99654 590620 135098
rect 590020 99418 590202 99654
rect 590438 99418 590620 99654
rect 590020 99334 590620 99418
rect 590020 99098 590202 99334
rect 590438 99098 590620 99334
rect 590020 63654 590620 99098
rect 590020 63418 590202 63654
rect 590438 63418 590620 63654
rect 590020 63334 590620 63418
rect 590020 63098 590202 63334
rect 590438 63098 590620 63334
rect 590020 27654 590620 63098
rect 590020 27418 590202 27654
rect 590438 27418 590620 27654
rect 590020 27334 590620 27418
rect 590020 27098 590202 27334
rect 590438 27098 590620 27334
rect 590020 -5046 590620 27098
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect 590960 697254 591560 709922
rect 590960 697018 591142 697254
rect 591378 697018 591560 697254
rect 590960 696934 591560 697018
rect 590960 696698 591142 696934
rect 591378 696698 591560 696934
rect 590960 661254 591560 696698
rect 590960 661018 591142 661254
rect 591378 661018 591560 661254
rect 590960 660934 591560 661018
rect 590960 660698 591142 660934
rect 591378 660698 591560 660934
rect 590960 625254 591560 660698
rect 590960 625018 591142 625254
rect 591378 625018 591560 625254
rect 590960 624934 591560 625018
rect 590960 624698 591142 624934
rect 591378 624698 591560 624934
rect 590960 589254 591560 624698
rect 590960 589018 591142 589254
rect 591378 589018 591560 589254
rect 590960 588934 591560 589018
rect 590960 588698 591142 588934
rect 591378 588698 591560 588934
rect 590960 553254 591560 588698
rect 590960 553018 591142 553254
rect 591378 553018 591560 553254
rect 590960 552934 591560 553018
rect 590960 552698 591142 552934
rect 591378 552698 591560 552934
rect 590960 517254 591560 552698
rect 590960 517018 591142 517254
rect 591378 517018 591560 517254
rect 590960 516934 591560 517018
rect 590960 516698 591142 516934
rect 591378 516698 591560 516934
rect 590960 481254 591560 516698
rect 590960 481018 591142 481254
rect 591378 481018 591560 481254
rect 590960 480934 591560 481018
rect 590960 480698 591142 480934
rect 591378 480698 591560 480934
rect 590960 445254 591560 480698
rect 590960 445018 591142 445254
rect 591378 445018 591560 445254
rect 590960 444934 591560 445018
rect 590960 444698 591142 444934
rect 591378 444698 591560 444934
rect 590960 409254 591560 444698
rect 590960 409018 591142 409254
rect 591378 409018 591560 409254
rect 590960 408934 591560 409018
rect 590960 408698 591142 408934
rect 591378 408698 591560 408934
rect 590960 373254 591560 408698
rect 590960 373018 591142 373254
rect 591378 373018 591560 373254
rect 590960 372934 591560 373018
rect 590960 372698 591142 372934
rect 591378 372698 591560 372934
rect 590960 337254 591560 372698
rect 590960 337018 591142 337254
rect 591378 337018 591560 337254
rect 590960 336934 591560 337018
rect 590960 336698 591142 336934
rect 591378 336698 591560 336934
rect 590960 301254 591560 336698
rect 590960 301018 591142 301254
rect 591378 301018 591560 301254
rect 590960 300934 591560 301018
rect 590960 300698 591142 300934
rect 591378 300698 591560 300934
rect 590960 265254 591560 300698
rect 590960 265018 591142 265254
rect 591378 265018 591560 265254
rect 590960 264934 591560 265018
rect 590960 264698 591142 264934
rect 591378 264698 591560 264934
rect 590960 229254 591560 264698
rect 590960 229018 591142 229254
rect 591378 229018 591560 229254
rect 590960 228934 591560 229018
rect 590960 228698 591142 228934
rect 591378 228698 591560 228934
rect 590960 193254 591560 228698
rect 590960 193018 591142 193254
rect 591378 193018 591560 193254
rect 590960 192934 591560 193018
rect 590960 192698 591142 192934
rect 591378 192698 591560 192934
rect 590960 157254 591560 192698
rect 590960 157018 591142 157254
rect 591378 157018 591560 157254
rect 590960 156934 591560 157018
rect 590960 156698 591142 156934
rect 591378 156698 591560 156934
rect 590960 121254 591560 156698
rect 590960 121018 591142 121254
rect 591378 121018 591560 121254
rect 590960 120934 591560 121018
rect 590960 120698 591142 120934
rect 591378 120698 591560 120934
rect 590960 85254 591560 120698
rect 590960 85018 591142 85254
rect 591378 85018 591560 85254
rect 590960 84934 591560 85018
rect 590960 84698 591142 84934
rect 591378 84698 591560 84934
rect 590960 49254 591560 84698
rect 590960 49018 591142 49254
rect 591378 49018 591560 49254
rect 590960 48934 591560 49018
rect 590960 48698 591142 48934
rect 591378 48698 591560 48934
rect 590960 13254 591560 48698
rect 590960 13018 591142 13254
rect 591378 13018 591560 13254
rect 590960 12934 591560 13018
rect 590960 12698 591142 12934
rect 591378 12698 591560 12934
rect 590960 -5986 591560 12698
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect 591900 679254 592500 710862
rect 591900 679018 592082 679254
rect 592318 679018 592500 679254
rect 591900 678934 592500 679018
rect 591900 678698 592082 678934
rect 592318 678698 592500 678934
rect 591900 643254 592500 678698
rect 591900 643018 592082 643254
rect 592318 643018 592500 643254
rect 591900 642934 592500 643018
rect 591900 642698 592082 642934
rect 592318 642698 592500 642934
rect 591900 607254 592500 642698
rect 591900 607018 592082 607254
rect 592318 607018 592500 607254
rect 591900 606934 592500 607018
rect 591900 606698 592082 606934
rect 592318 606698 592500 606934
rect 591900 571254 592500 606698
rect 591900 571018 592082 571254
rect 592318 571018 592500 571254
rect 591900 570934 592500 571018
rect 591900 570698 592082 570934
rect 592318 570698 592500 570934
rect 591900 535254 592500 570698
rect 591900 535018 592082 535254
rect 592318 535018 592500 535254
rect 591900 534934 592500 535018
rect 591900 534698 592082 534934
rect 592318 534698 592500 534934
rect 591900 499254 592500 534698
rect 591900 499018 592082 499254
rect 592318 499018 592500 499254
rect 591900 498934 592500 499018
rect 591900 498698 592082 498934
rect 592318 498698 592500 498934
rect 591900 463254 592500 498698
rect 591900 463018 592082 463254
rect 592318 463018 592500 463254
rect 591900 462934 592500 463018
rect 591900 462698 592082 462934
rect 592318 462698 592500 462934
rect 591900 427254 592500 462698
rect 591900 427018 592082 427254
rect 592318 427018 592500 427254
rect 591900 426934 592500 427018
rect 591900 426698 592082 426934
rect 592318 426698 592500 426934
rect 591900 391254 592500 426698
rect 591900 391018 592082 391254
rect 592318 391018 592500 391254
rect 591900 390934 592500 391018
rect 591900 390698 592082 390934
rect 592318 390698 592500 390934
rect 591900 355254 592500 390698
rect 591900 355018 592082 355254
rect 592318 355018 592500 355254
rect 591900 354934 592500 355018
rect 591900 354698 592082 354934
rect 592318 354698 592500 354934
rect 591900 319254 592500 354698
rect 591900 319018 592082 319254
rect 592318 319018 592500 319254
rect 591900 318934 592500 319018
rect 591900 318698 592082 318934
rect 592318 318698 592500 318934
rect 591900 283254 592500 318698
rect 591900 283018 592082 283254
rect 592318 283018 592500 283254
rect 591900 282934 592500 283018
rect 591900 282698 592082 282934
rect 592318 282698 592500 282934
rect 591900 247254 592500 282698
rect 591900 247018 592082 247254
rect 592318 247018 592500 247254
rect 591900 246934 592500 247018
rect 591900 246698 592082 246934
rect 592318 246698 592500 246934
rect 591900 211254 592500 246698
rect 591900 211018 592082 211254
rect 592318 211018 592500 211254
rect 591900 210934 592500 211018
rect 591900 210698 592082 210934
rect 592318 210698 592500 210934
rect 591900 175254 592500 210698
rect 591900 175018 592082 175254
rect 592318 175018 592500 175254
rect 591900 174934 592500 175018
rect 591900 174698 592082 174934
rect 592318 174698 592500 174934
rect 591900 139254 592500 174698
rect 591900 139018 592082 139254
rect 592318 139018 592500 139254
rect 591900 138934 592500 139018
rect 591900 138698 592082 138934
rect 592318 138698 592500 138934
rect 591900 103254 592500 138698
rect 591900 103018 592082 103254
rect 592318 103018 592500 103254
rect 591900 102934 592500 103018
rect 591900 102698 592082 102934
rect 592318 102698 592500 102934
rect 591900 67254 592500 102698
rect 591900 67018 592082 67254
rect 592318 67018 592500 67254
rect 591900 66934 592500 67018
rect 591900 66698 592082 66934
rect 592318 66698 592500 66934
rect 591900 31254 592500 66698
rect 591900 31018 592082 31254
rect 592318 31018 592500 31254
rect 591900 30934 592500 31018
rect 591900 30698 592082 30934
rect 592318 30698 592500 30934
rect 569604 -7162 569786 -6926
rect 570022 -7162 570204 -6926
rect 569604 -7246 570204 -7162
rect 569604 -7482 569786 -7246
rect 570022 -7482 570204 -7246
rect 569604 -7504 570204 -7482
rect 591900 -6926 592500 30698
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect -8394 679018 -8158 679254
rect -8394 678698 -8158 678934
rect -8394 643018 -8158 643254
rect -8394 642698 -8158 642934
rect -8394 607018 -8158 607254
rect -8394 606698 -8158 606934
rect -8394 571018 -8158 571254
rect -8394 570698 -8158 570934
rect -8394 535018 -8158 535254
rect -8394 534698 -8158 534934
rect -8394 499018 -8158 499254
rect -8394 498698 -8158 498934
rect -8394 463018 -8158 463254
rect -8394 462698 -8158 462934
rect -8394 427018 -8158 427254
rect -8394 426698 -8158 426934
rect -8394 391018 -8158 391254
rect -8394 390698 -8158 390934
rect -8394 355018 -8158 355254
rect -8394 354698 -8158 354934
rect -8394 319018 -8158 319254
rect -8394 318698 -8158 318934
rect -8394 283018 -8158 283254
rect -8394 282698 -8158 282934
rect -8394 247018 -8158 247254
rect -8394 246698 -8158 246934
rect -8394 211018 -8158 211254
rect -8394 210698 -8158 210934
rect -8394 175018 -8158 175254
rect -8394 174698 -8158 174934
rect -8394 139018 -8158 139254
rect -8394 138698 -8158 138934
rect -8394 103018 -8158 103254
rect -8394 102698 -8158 102934
rect -8394 67018 -8158 67254
rect -8394 66698 -8158 66934
rect -8394 31018 -8158 31254
rect -8394 30698 -8158 30934
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 11786 710242 12022 710478
rect 11786 709922 12022 710158
rect -7454 697018 -7218 697254
rect -7454 696698 -7218 696934
rect -7454 661018 -7218 661254
rect -7454 660698 -7218 660934
rect -7454 625018 -7218 625254
rect -7454 624698 -7218 624934
rect -7454 589018 -7218 589254
rect -7454 588698 -7218 588934
rect -7454 553018 -7218 553254
rect -7454 552698 -7218 552934
rect -7454 517018 -7218 517254
rect -7454 516698 -7218 516934
rect -7454 481018 -7218 481254
rect -7454 480698 -7218 480934
rect -7454 445018 -7218 445254
rect -7454 444698 -7218 444934
rect -7454 409018 -7218 409254
rect -7454 408698 -7218 408934
rect -7454 373018 -7218 373254
rect -7454 372698 -7218 372934
rect -7454 337018 -7218 337254
rect -7454 336698 -7218 336934
rect -7454 301018 -7218 301254
rect -7454 300698 -7218 300934
rect -7454 265018 -7218 265254
rect -7454 264698 -7218 264934
rect -7454 229018 -7218 229254
rect -7454 228698 -7218 228934
rect -7454 193018 -7218 193254
rect -7454 192698 -7218 192934
rect -7454 157018 -7218 157254
rect -7454 156698 -7218 156934
rect -7454 121018 -7218 121254
rect -7454 120698 -7218 120934
rect -7454 85018 -7218 85254
rect -7454 84698 -7218 84934
rect -7454 49018 -7218 49254
rect -7454 48698 -7218 48934
rect -7454 13018 -7218 13254
rect -7454 12698 -7218 12934
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect -6514 675418 -6278 675654
rect -6514 675098 -6278 675334
rect -6514 639418 -6278 639654
rect -6514 639098 -6278 639334
rect -6514 603418 -6278 603654
rect -6514 603098 -6278 603334
rect -6514 567418 -6278 567654
rect -6514 567098 -6278 567334
rect -6514 531418 -6278 531654
rect -6514 531098 -6278 531334
rect -6514 495418 -6278 495654
rect -6514 495098 -6278 495334
rect -6514 459418 -6278 459654
rect -6514 459098 -6278 459334
rect -6514 423418 -6278 423654
rect -6514 423098 -6278 423334
rect -6514 387418 -6278 387654
rect -6514 387098 -6278 387334
rect -6514 351418 -6278 351654
rect -6514 351098 -6278 351334
rect -6514 315418 -6278 315654
rect -6514 315098 -6278 315334
rect -6514 279418 -6278 279654
rect -6514 279098 -6278 279334
rect -6514 243418 -6278 243654
rect -6514 243098 -6278 243334
rect -6514 207418 -6278 207654
rect -6514 207098 -6278 207334
rect -6514 171418 -6278 171654
rect -6514 171098 -6278 171334
rect -6514 135418 -6278 135654
rect -6514 135098 -6278 135334
rect -6514 99418 -6278 99654
rect -6514 99098 -6278 99334
rect -6514 63418 -6278 63654
rect -6514 63098 -6278 63334
rect -6514 27418 -6278 27654
rect -6514 27098 -6278 27334
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 8186 708362 8422 708598
rect 8186 708042 8422 708278
rect -5574 693418 -5338 693654
rect -5574 693098 -5338 693334
rect -5574 657418 -5338 657654
rect -5574 657098 -5338 657334
rect -5574 621418 -5338 621654
rect -5574 621098 -5338 621334
rect -5574 585418 -5338 585654
rect -5574 585098 -5338 585334
rect -5574 549418 -5338 549654
rect -5574 549098 -5338 549334
rect -5574 513418 -5338 513654
rect -5574 513098 -5338 513334
rect -5574 477418 -5338 477654
rect -5574 477098 -5338 477334
rect -5574 441418 -5338 441654
rect -5574 441098 -5338 441334
rect -5574 405418 -5338 405654
rect -5574 405098 -5338 405334
rect -5574 369418 -5338 369654
rect -5574 369098 -5338 369334
rect -5574 333418 -5338 333654
rect -5574 333098 -5338 333334
rect -5574 297418 -5338 297654
rect -5574 297098 -5338 297334
rect -5574 261418 -5338 261654
rect -5574 261098 -5338 261334
rect -5574 225418 -5338 225654
rect -5574 225098 -5338 225334
rect -5574 189418 -5338 189654
rect -5574 189098 -5338 189334
rect -5574 153418 -5338 153654
rect -5574 153098 -5338 153334
rect -5574 117418 -5338 117654
rect -5574 117098 -5338 117334
rect -5574 81418 -5338 81654
rect -5574 81098 -5338 81334
rect -5574 45418 -5338 45654
rect -5574 45098 -5338 45334
rect -5574 9418 -5338 9654
rect -5574 9098 -5338 9334
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect -4634 671818 -4398 672054
rect -4634 671498 -4398 671734
rect -4634 635818 -4398 636054
rect -4634 635498 -4398 635734
rect -4634 599818 -4398 600054
rect -4634 599498 -4398 599734
rect -4634 563818 -4398 564054
rect -4634 563498 -4398 563734
rect -4634 527818 -4398 528054
rect -4634 527498 -4398 527734
rect -4634 491818 -4398 492054
rect -4634 491498 -4398 491734
rect -4634 455818 -4398 456054
rect -4634 455498 -4398 455734
rect -4634 419818 -4398 420054
rect -4634 419498 -4398 419734
rect -4634 383818 -4398 384054
rect -4634 383498 -4398 383734
rect -4634 347818 -4398 348054
rect -4634 347498 -4398 347734
rect -4634 311818 -4398 312054
rect -4634 311498 -4398 311734
rect -4634 275818 -4398 276054
rect -4634 275498 -4398 275734
rect -4634 239818 -4398 240054
rect -4634 239498 -4398 239734
rect -4634 203818 -4398 204054
rect -4634 203498 -4398 203734
rect -4634 167818 -4398 168054
rect -4634 167498 -4398 167734
rect -4634 131818 -4398 132054
rect -4634 131498 -4398 131734
rect -4634 95818 -4398 96054
rect -4634 95498 -4398 95734
rect -4634 59818 -4398 60054
rect -4634 59498 -4398 59734
rect -4634 23818 -4398 24054
rect -4634 23498 -4398 23734
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 4586 706482 4822 706718
rect 4586 706162 4822 706398
rect -3694 689818 -3458 690054
rect -3694 689498 -3458 689734
rect -3694 653818 -3458 654054
rect -3694 653498 -3458 653734
rect -3694 617818 -3458 618054
rect -3694 617498 -3458 617734
rect -3694 581818 -3458 582054
rect -3694 581498 -3458 581734
rect -3694 545818 -3458 546054
rect -3694 545498 -3458 545734
rect -3694 509818 -3458 510054
rect -3694 509498 -3458 509734
rect -3694 473818 -3458 474054
rect -3694 473498 -3458 473734
rect -3694 437818 -3458 438054
rect -3694 437498 -3458 437734
rect -3694 401818 -3458 402054
rect -3694 401498 -3458 401734
rect -3694 365818 -3458 366054
rect -3694 365498 -3458 365734
rect -3694 329818 -3458 330054
rect -3694 329498 -3458 329734
rect -3694 293818 -3458 294054
rect -3694 293498 -3458 293734
rect -3694 257818 -3458 258054
rect -3694 257498 -3458 257734
rect -3694 221818 -3458 222054
rect -3694 221498 -3458 221734
rect -3694 185818 -3458 186054
rect -3694 185498 -3458 185734
rect -3694 149818 -3458 150054
rect -3694 149498 -3458 149734
rect -3694 113818 -3458 114054
rect -3694 113498 -3458 113734
rect -3694 77818 -3458 78054
rect -3694 77498 -3458 77734
rect -3694 41818 -3458 42054
rect -3694 41498 -3458 41734
rect -3694 5818 -3458 6054
rect -3694 5498 -3458 5734
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 29786 711182 30022 711418
rect 29786 710862 30022 711098
rect 26186 709302 26422 709538
rect 26186 708982 26422 709218
rect 22586 707422 22822 707658
rect 22586 707102 22822 707338
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 47786 710242 48022 710478
rect 47786 709922 48022 710158
rect 44186 708362 44422 708598
rect 44186 708042 44422 708278
rect 40586 706482 40822 706718
rect 40586 706162 40822 706398
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect 65786 711182 66022 711418
rect 65786 710862 66022 711098
rect 62186 709302 62422 709538
rect 62186 708982 62422 709218
rect 58586 707422 58822 707658
rect 58586 707102 58822 707338
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 83786 710242 84022 710478
rect 83786 709922 84022 710158
rect 80186 708362 80422 708598
rect 80186 708042 80422 708278
rect 76586 706482 76822 706718
rect 76586 706162 76822 706398
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 101786 711182 102022 711418
rect 101786 710862 102022 711098
rect 98186 709302 98422 709538
rect 98186 708982 98422 709218
rect 94586 707422 94822 707658
rect 94586 707102 94822 707338
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 119786 710242 120022 710478
rect 119786 709922 120022 710158
rect 116186 708362 116422 708598
rect 116186 708042 116422 708278
rect 112586 706482 112822 706718
rect 112586 706162 112822 706398
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 137786 711182 138022 711418
rect 137786 710862 138022 711098
rect 134186 709302 134422 709538
rect 134186 708982 134422 709218
rect 130586 707422 130822 707658
rect 130586 707102 130822 707338
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 155786 710242 156022 710478
rect 155786 709922 156022 710158
rect 152186 708362 152422 708598
rect 152186 708042 152422 708278
rect 148586 706482 148822 706718
rect 148586 706162 148822 706398
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 173786 711182 174022 711418
rect 173786 710862 174022 711098
rect 170186 709302 170422 709538
rect 170186 708982 170422 709218
rect 166586 707422 166822 707658
rect 166586 707102 166822 707338
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 191786 710242 192022 710478
rect 191786 709922 192022 710158
rect 188186 708362 188422 708598
rect 188186 708042 188422 708278
rect 184586 706482 184822 706718
rect 184586 706162 184822 706398
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 209786 711182 210022 711418
rect 209786 710862 210022 711098
rect 206186 709302 206422 709538
rect 206186 708982 206422 709218
rect 202586 707422 202822 707658
rect 202586 707102 202822 707338
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 227786 710242 228022 710478
rect 227786 709922 228022 710158
rect 224186 708362 224422 708598
rect 224186 708042 224422 708278
rect 220586 706482 220822 706718
rect 220586 706162 220822 706398
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 245786 711182 246022 711418
rect 245786 710862 246022 711098
rect 242186 709302 242422 709538
rect 242186 708982 242422 709218
rect 238586 707422 238822 707658
rect 238586 707102 238822 707338
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 263786 710242 264022 710478
rect 263786 709922 264022 710158
rect 260186 708362 260422 708598
rect 260186 708042 260422 708278
rect 256586 706482 256822 706718
rect 256586 706162 256822 706398
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 281786 711182 282022 711418
rect 281786 710862 282022 711098
rect 278186 709302 278422 709538
rect 278186 708982 278422 709218
rect 274586 707422 274822 707658
rect 274586 707102 274822 707338
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 299786 710242 300022 710478
rect 299786 709922 300022 710158
rect 296186 708362 296422 708598
rect 296186 708042 296422 708278
rect 292586 706482 292822 706718
rect 292586 706162 292822 706398
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 317786 711182 318022 711418
rect 317786 710862 318022 711098
rect 314186 709302 314422 709538
rect 314186 708982 314422 709218
rect 310586 707422 310822 707658
rect 310586 707102 310822 707338
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 335786 710242 336022 710478
rect 335786 709922 336022 710158
rect 332186 708362 332422 708598
rect 332186 708042 332422 708278
rect 328586 706482 328822 706718
rect 328586 706162 328822 706398
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 353786 711182 354022 711418
rect 353786 710862 354022 711098
rect 350186 709302 350422 709538
rect 350186 708982 350422 709218
rect 346586 707422 346822 707658
rect 346586 707102 346822 707338
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 371786 710242 372022 710478
rect 371786 709922 372022 710158
rect 368186 708362 368422 708598
rect 368186 708042 368422 708278
rect 364586 706482 364822 706718
rect 364586 706162 364822 706398
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 389786 711182 390022 711418
rect 389786 710862 390022 711098
rect 386186 709302 386422 709538
rect 386186 708982 386422 709218
rect 382586 707422 382822 707658
rect 382586 707102 382822 707338
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 407786 710242 408022 710478
rect 407786 709922 408022 710158
rect 404186 708362 404422 708598
rect 404186 708042 404422 708278
rect 400586 706482 400822 706718
rect 400586 706162 400822 706398
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 425786 711182 426022 711418
rect 425786 710862 426022 711098
rect 422186 709302 422422 709538
rect 422186 708982 422422 709218
rect 418586 707422 418822 707658
rect 418586 707102 418822 707338
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 443786 710242 444022 710478
rect 443786 709922 444022 710158
rect 440186 708362 440422 708598
rect 440186 708042 440422 708278
rect 436586 706482 436822 706718
rect 436586 706162 436822 706398
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 461786 711182 462022 711418
rect 461786 710862 462022 711098
rect 458186 709302 458422 709538
rect 458186 708982 458422 709218
rect 454586 707422 454822 707658
rect 454586 707102 454822 707338
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 479786 710242 480022 710478
rect 479786 709922 480022 710158
rect 476186 708362 476422 708598
rect 476186 708042 476422 708278
rect 472586 706482 472822 706718
rect 472586 706162 472822 706398
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 497786 711182 498022 711418
rect 497786 710862 498022 711098
rect 494186 709302 494422 709538
rect 494186 708982 494422 709218
rect 490586 707422 490822 707658
rect 490586 707102 490822 707338
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 515786 710242 516022 710478
rect 515786 709922 516022 710158
rect 512186 708362 512422 708598
rect 512186 708042 512422 708278
rect 508586 706482 508822 706718
rect 508586 706162 508822 706398
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 533786 711182 534022 711418
rect 533786 710862 534022 711098
rect 530186 709302 530422 709538
rect 530186 708982 530422 709218
rect 526586 707422 526822 707658
rect 526586 707102 526822 707338
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 551786 710242 552022 710478
rect 551786 709922 552022 710158
rect 548186 708362 548422 708598
rect 548186 708042 548422 708278
rect 544586 706482 544822 706718
rect 544586 706162 544822 706398
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 569786 711182 570022 711418
rect 569786 710862 570022 711098
rect 566186 709302 566422 709538
rect 566186 708982 566422 709218
rect 562586 707422 562822 707658
rect 562586 707102 562822 707338
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 580586 706482 580822 706718
rect 580586 706162 580822 706398
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 35506 596218 35742 596454
rect 35506 595898 35742 596134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 545562 632214 545798 632450
rect 545562 631894 545798 632130
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect 545990 578216 546226 578452
rect 545990 577896 546226 578132
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect 34600 470218 34836 470454
rect 34600 469898 34836 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect 35034 416220 35270 416456
rect 35034 415900 35270 416136
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 545560 416210 545796 416446
rect 545560 415890 545796 416126
rect 545956 398224 546192 398460
rect 545956 397904 546192 398140
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 544412 236222 544648 236458
rect 544412 235902 544648 236138
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect 544876 182232 545112 182468
rect 544876 181912 545112 182148
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 4586 -2462 4822 -2226
rect 4586 -2782 4822 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 8186 -4342 8422 -4106
rect 8186 -4662 8422 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 22586 -3402 22822 -3166
rect 22586 -3722 22822 -3486
rect 26186 -5282 26422 -5046
rect 26186 -5602 26422 -5366
rect 11786 -6222 12022 -5986
rect 11786 -6542 12022 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 -2462 40822 -2226
rect 40586 -2782 40822 -2546
rect 44186 -4342 44422 -4106
rect 44186 -4662 44422 -4426
rect 29786 -7162 30022 -6926
rect 29786 -7482 30022 -7246
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 58586 -3402 58822 -3166
rect 58586 -3722 58822 -3486
rect 62186 -5282 62422 -5046
rect 62186 -5602 62422 -5366
rect 47786 -6222 48022 -5986
rect 47786 -6542 48022 -6306
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 -2462 76822 -2226
rect 76586 -2782 76822 -2546
rect 80186 -4342 80422 -4106
rect 80186 -4662 80422 -4426
rect 65786 -7162 66022 -6926
rect 65786 -7482 66022 -7246
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 94586 -3402 94822 -3166
rect 94586 -3722 94822 -3486
rect 98186 -5282 98422 -5046
rect 98186 -5602 98422 -5366
rect 83786 -6222 84022 -5986
rect 83786 -6542 84022 -6306
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 -2462 112822 -2226
rect 112586 -2782 112822 -2546
rect 116186 -4342 116422 -4106
rect 116186 -4662 116422 -4426
rect 101786 -7162 102022 -6926
rect 101786 -7482 102022 -7246
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 130586 -3402 130822 -3166
rect 130586 -3722 130822 -3486
rect 134186 -5282 134422 -5046
rect 134186 -5602 134422 -5366
rect 119786 -6222 120022 -5986
rect 119786 -6542 120022 -6306
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 -2462 148822 -2226
rect 148586 -2782 148822 -2546
rect 152186 -4342 152422 -4106
rect 152186 -4662 152422 -4426
rect 137786 -7162 138022 -6926
rect 137786 -7482 138022 -7246
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 166586 -3402 166822 -3166
rect 166586 -3722 166822 -3486
rect 170186 -5282 170422 -5046
rect 170186 -5602 170422 -5366
rect 155786 -6222 156022 -5986
rect 155786 -6542 156022 -6306
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 -2462 184822 -2226
rect 184586 -2782 184822 -2546
rect 188186 -4342 188422 -4106
rect 188186 -4662 188422 -4426
rect 173786 -7162 174022 -6926
rect 173786 -7482 174022 -7246
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 202586 -3402 202822 -3166
rect 202586 -3722 202822 -3486
rect 206186 -5282 206422 -5046
rect 206186 -5602 206422 -5366
rect 191786 -6222 192022 -5986
rect 191786 -6542 192022 -6306
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 -2462 220822 -2226
rect 220586 -2782 220822 -2546
rect 224186 -4342 224422 -4106
rect 224186 -4662 224422 -4426
rect 209786 -7162 210022 -6926
rect 209786 -7482 210022 -7246
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 238586 -3402 238822 -3166
rect 238586 -3722 238822 -3486
rect 242186 -5282 242422 -5046
rect 242186 -5602 242422 -5366
rect 227786 -6222 228022 -5986
rect 227786 -6542 228022 -6306
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 -2462 256822 -2226
rect 256586 -2782 256822 -2546
rect 260186 -4342 260422 -4106
rect 260186 -4662 260422 -4426
rect 245786 -7162 246022 -6926
rect 245786 -7482 246022 -7246
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 274586 -3402 274822 -3166
rect 274586 -3722 274822 -3486
rect 278186 -5282 278422 -5046
rect 278186 -5602 278422 -5366
rect 263786 -6222 264022 -5986
rect 263786 -6542 264022 -6306
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 -2462 292822 -2226
rect 292586 -2782 292822 -2546
rect 296186 -4342 296422 -4106
rect 296186 -4662 296422 -4426
rect 281786 -7162 282022 -6926
rect 281786 -7482 282022 -7246
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 310586 -3402 310822 -3166
rect 310586 -3722 310822 -3486
rect 314186 -5282 314422 -5046
rect 314186 -5602 314422 -5366
rect 299786 -6222 300022 -5986
rect 299786 -6542 300022 -6306
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 -2462 328822 -2226
rect 328586 -2782 328822 -2546
rect 332186 -4342 332422 -4106
rect 332186 -4662 332422 -4426
rect 317786 -7162 318022 -6926
rect 317786 -7482 318022 -7246
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 346586 -3402 346822 -3166
rect 346586 -3722 346822 -3486
rect 350186 -5282 350422 -5046
rect 350186 -5602 350422 -5366
rect 335786 -6222 336022 -5986
rect 335786 -6542 336022 -6306
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 -2462 364822 -2226
rect 364586 -2782 364822 -2546
rect 368186 -4342 368422 -4106
rect 368186 -4662 368422 -4426
rect 353786 -7162 354022 -6926
rect 353786 -7482 354022 -7246
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 382586 -3402 382822 -3166
rect 382586 -3722 382822 -3486
rect 386186 -5282 386422 -5046
rect 386186 -5602 386422 -5366
rect 371786 -6222 372022 -5986
rect 371786 -6542 372022 -6306
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 -2462 400822 -2226
rect 400586 -2782 400822 -2546
rect 404186 -4342 404422 -4106
rect 404186 -4662 404422 -4426
rect 389786 -7162 390022 -6926
rect 389786 -7482 390022 -7246
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 418586 -3402 418822 -3166
rect 418586 -3722 418822 -3486
rect 422186 -5282 422422 -5046
rect 422186 -5602 422422 -5366
rect 407786 -6222 408022 -5986
rect 407786 -6542 408022 -6306
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 -2462 436822 -2226
rect 436586 -2782 436822 -2546
rect 440186 -4342 440422 -4106
rect 440186 -4662 440422 -4426
rect 425786 -7162 426022 -6926
rect 425786 -7482 426022 -7246
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 454586 -3402 454822 -3166
rect 454586 -3722 454822 -3486
rect 458186 -5282 458422 -5046
rect 458186 -5602 458422 -5366
rect 443786 -6222 444022 -5986
rect 443786 -6542 444022 -6306
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 -2462 472822 -2226
rect 472586 -2782 472822 -2546
rect 476186 -4342 476422 -4106
rect 476186 -4662 476422 -4426
rect 461786 -7162 462022 -6926
rect 461786 -7482 462022 -7246
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 490586 -3402 490822 -3166
rect 490586 -3722 490822 -3486
rect 494186 -5282 494422 -5046
rect 494186 -5602 494422 -5366
rect 479786 -6222 480022 -5986
rect 479786 -6542 480022 -6306
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 -2462 508822 -2226
rect 508586 -2782 508822 -2546
rect 512186 -4342 512422 -4106
rect 512186 -4662 512422 -4426
rect 497786 -7162 498022 -6926
rect 497786 -7482 498022 -7246
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 526586 -3402 526822 -3166
rect 526586 -3722 526822 -3486
rect 530186 -5282 530422 -5046
rect 530186 -5602 530422 -5366
rect 515786 -6222 516022 -5986
rect 515786 -6542 516022 -6306
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 -2462 544822 -2226
rect 544586 -2782 544822 -2546
rect 548186 -4342 548422 -4106
rect 548186 -4662 548422 -4426
rect 533786 -7162 534022 -6926
rect 533786 -7482 534022 -7246
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 562586 -3402 562822 -3166
rect 562586 -3722 562822 -3486
rect 566186 -5282 566422 -5046
rect 566186 -5602 566422 -5366
rect 551786 -6222 552022 -5986
rect 551786 -6542 552022 -6306
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 587382 689818 587618 690054
rect 587382 689498 587618 689734
rect 587382 653818 587618 654054
rect 587382 653498 587618 653734
rect 587382 617818 587618 618054
rect 587382 617498 587618 617734
rect 587382 581818 587618 582054
rect 587382 581498 587618 581734
rect 587382 545818 587618 546054
rect 587382 545498 587618 545734
rect 587382 509818 587618 510054
rect 587382 509498 587618 509734
rect 587382 473818 587618 474054
rect 587382 473498 587618 473734
rect 587382 437818 587618 438054
rect 587382 437498 587618 437734
rect 587382 401818 587618 402054
rect 587382 401498 587618 401734
rect 587382 365818 587618 366054
rect 587382 365498 587618 365734
rect 587382 329818 587618 330054
rect 587382 329498 587618 329734
rect 587382 293818 587618 294054
rect 587382 293498 587618 293734
rect 587382 257818 587618 258054
rect 587382 257498 587618 257734
rect 587382 221818 587618 222054
rect 587382 221498 587618 221734
rect 587382 185818 587618 186054
rect 587382 185498 587618 185734
rect 587382 149818 587618 150054
rect 587382 149498 587618 149734
rect 587382 113818 587618 114054
rect 587382 113498 587618 113734
rect 587382 77818 587618 78054
rect 587382 77498 587618 77734
rect 587382 41818 587618 42054
rect 587382 41498 587618 41734
rect 587382 5818 587618 6054
rect 587382 5498 587618 5734
rect 580586 -2462 580822 -2226
rect 580586 -2782 580822 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 671818 588558 672054
rect 588322 671498 588558 671734
rect 588322 635818 588558 636054
rect 588322 635498 588558 635734
rect 588322 599818 588558 600054
rect 588322 599498 588558 599734
rect 588322 563818 588558 564054
rect 588322 563498 588558 563734
rect 588322 527818 588558 528054
rect 588322 527498 588558 527734
rect 588322 491818 588558 492054
rect 588322 491498 588558 491734
rect 588322 455818 588558 456054
rect 588322 455498 588558 455734
rect 588322 419818 588558 420054
rect 588322 419498 588558 419734
rect 588322 383818 588558 384054
rect 588322 383498 588558 383734
rect 588322 347818 588558 348054
rect 588322 347498 588558 347734
rect 588322 311818 588558 312054
rect 588322 311498 588558 311734
rect 588322 275818 588558 276054
rect 588322 275498 588558 275734
rect 588322 239818 588558 240054
rect 588322 239498 588558 239734
rect 588322 203818 588558 204054
rect 588322 203498 588558 203734
rect 588322 167818 588558 168054
rect 588322 167498 588558 167734
rect 588322 131818 588558 132054
rect 588322 131498 588558 131734
rect 588322 95818 588558 96054
rect 588322 95498 588558 95734
rect 588322 59818 588558 60054
rect 588322 59498 588558 59734
rect 588322 23818 588558 24054
rect 588322 23498 588558 23734
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect 589262 693418 589498 693654
rect 589262 693098 589498 693334
rect 589262 657418 589498 657654
rect 589262 657098 589498 657334
rect 589262 621418 589498 621654
rect 589262 621098 589498 621334
rect 589262 585418 589498 585654
rect 589262 585098 589498 585334
rect 589262 549418 589498 549654
rect 589262 549098 589498 549334
rect 589262 513418 589498 513654
rect 589262 513098 589498 513334
rect 589262 477418 589498 477654
rect 589262 477098 589498 477334
rect 589262 441418 589498 441654
rect 589262 441098 589498 441334
rect 589262 405418 589498 405654
rect 589262 405098 589498 405334
rect 589262 369418 589498 369654
rect 589262 369098 589498 369334
rect 589262 333418 589498 333654
rect 589262 333098 589498 333334
rect 589262 297418 589498 297654
rect 589262 297098 589498 297334
rect 589262 261418 589498 261654
rect 589262 261098 589498 261334
rect 589262 225418 589498 225654
rect 589262 225098 589498 225334
rect 589262 189418 589498 189654
rect 589262 189098 589498 189334
rect 589262 153418 589498 153654
rect 589262 153098 589498 153334
rect 589262 117418 589498 117654
rect 589262 117098 589498 117334
rect 589262 81418 589498 81654
rect 589262 81098 589498 81334
rect 589262 45418 589498 45654
rect 589262 45098 589498 45334
rect 589262 9418 589498 9654
rect 589262 9098 589498 9334
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect 590202 675418 590438 675654
rect 590202 675098 590438 675334
rect 590202 639418 590438 639654
rect 590202 639098 590438 639334
rect 590202 603418 590438 603654
rect 590202 603098 590438 603334
rect 590202 567418 590438 567654
rect 590202 567098 590438 567334
rect 590202 531418 590438 531654
rect 590202 531098 590438 531334
rect 590202 495418 590438 495654
rect 590202 495098 590438 495334
rect 590202 459418 590438 459654
rect 590202 459098 590438 459334
rect 590202 423418 590438 423654
rect 590202 423098 590438 423334
rect 590202 387418 590438 387654
rect 590202 387098 590438 387334
rect 590202 351418 590438 351654
rect 590202 351098 590438 351334
rect 590202 315418 590438 315654
rect 590202 315098 590438 315334
rect 590202 279418 590438 279654
rect 590202 279098 590438 279334
rect 590202 243418 590438 243654
rect 590202 243098 590438 243334
rect 590202 207418 590438 207654
rect 590202 207098 590438 207334
rect 590202 171418 590438 171654
rect 590202 171098 590438 171334
rect 590202 135418 590438 135654
rect 590202 135098 590438 135334
rect 590202 99418 590438 99654
rect 590202 99098 590438 99334
rect 590202 63418 590438 63654
rect 590202 63098 590438 63334
rect 590202 27418 590438 27654
rect 590202 27098 590438 27334
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect 591142 697018 591378 697254
rect 591142 696698 591378 696934
rect 591142 661018 591378 661254
rect 591142 660698 591378 660934
rect 591142 625018 591378 625254
rect 591142 624698 591378 624934
rect 591142 589018 591378 589254
rect 591142 588698 591378 588934
rect 591142 553018 591378 553254
rect 591142 552698 591378 552934
rect 591142 517018 591378 517254
rect 591142 516698 591378 516934
rect 591142 481018 591378 481254
rect 591142 480698 591378 480934
rect 591142 445018 591378 445254
rect 591142 444698 591378 444934
rect 591142 409018 591378 409254
rect 591142 408698 591378 408934
rect 591142 373018 591378 373254
rect 591142 372698 591378 372934
rect 591142 337018 591378 337254
rect 591142 336698 591378 336934
rect 591142 301018 591378 301254
rect 591142 300698 591378 300934
rect 591142 265018 591378 265254
rect 591142 264698 591378 264934
rect 591142 229018 591378 229254
rect 591142 228698 591378 228934
rect 591142 193018 591378 193254
rect 591142 192698 591378 192934
rect 591142 157018 591378 157254
rect 591142 156698 591378 156934
rect 591142 121018 591378 121254
rect 591142 120698 591378 120934
rect 591142 85018 591378 85254
rect 591142 84698 591378 84934
rect 591142 49018 591378 49254
rect 591142 48698 591378 48934
rect 591142 13018 591378 13254
rect 591142 12698 591378 12934
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect 592082 679018 592318 679254
rect 592082 678698 592318 678934
rect 592082 643018 592318 643254
rect 592082 642698 592318 642934
rect 592082 607018 592318 607254
rect 592082 606698 592318 606934
rect 592082 571018 592318 571254
rect 592082 570698 592318 570934
rect 592082 535018 592318 535254
rect 592082 534698 592318 534934
rect 592082 499018 592318 499254
rect 592082 498698 592318 498934
rect 592082 463018 592318 463254
rect 592082 462698 592318 462934
rect 592082 427018 592318 427254
rect 592082 426698 592318 426934
rect 592082 391018 592318 391254
rect 592082 390698 592318 390934
rect 592082 355018 592318 355254
rect 592082 354698 592318 354934
rect 592082 319018 592318 319254
rect 592082 318698 592318 318934
rect 592082 283018 592318 283254
rect 592082 282698 592318 282934
rect 592082 247018 592318 247254
rect 592082 246698 592318 246934
rect 592082 211018 592318 211254
rect 592082 210698 592318 210934
rect 592082 175018 592318 175254
rect 592082 174698 592318 174934
rect 592082 139018 592318 139254
rect 592082 138698 592318 138934
rect 592082 103018 592318 103254
rect 592082 102698 592318 102934
rect 592082 67018 592318 67254
rect 592082 66698 592318 66934
rect 592082 31018 592318 31254
rect 592082 30698 592318 30934
rect 569786 -7162 570022 -6926
rect 569786 -7482 570022 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 29604 711440 30204 711442
rect 65604 711440 66204 711442
rect 101604 711440 102204 711442
rect 137604 711440 138204 711442
rect 173604 711440 174204 711442
rect 209604 711440 210204 711442
rect 245604 711440 246204 711442
rect 281604 711440 282204 711442
rect 317604 711440 318204 711442
rect 353604 711440 354204 711442
rect 389604 711440 390204 711442
rect 425604 711440 426204 711442
rect 461604 711440 462204 711442
rect 497604 711440 498204 711442
rect 533604 711440 534204 711442
rect 569604 711440 570204 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 29786 711418
rect 30022 711182 65786 711418
rect 66022 711182 101786 711418
rect 102022 711182 137786 711418
rect 138022 711182 173786 711418
rect 174022 711182 209786 711418
rect 210022 711182 245786 711418
rect 246022 711182 281786 711418
rect 282022 711182 317786 711418
rect 318022 711182 353786 711418
rect 354022 711182 389786 711418
rect 390022 711182 425786 711418
rect 426022 711182 461786 711418
rect 462022 711182 497786 711418
rect 498022 711182 533786 711418
rect 534022 711182 569786 711418
rect 570022 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 29786 711098
rect 30022 710862 65786 711098
rect 66022 710862 101786 711098
rect 102022 710862 137786 711098
rect 138022 710862 173786 711098
rect 174022 710862 209786 711098
rect 210022 710862 245786 711098
rect 246022 710862 281786 711098
rect 282022 710862 317786 711098
rect 318022 710862 353786 711098
rect 354022 710862 389786 711098
rect 390022 710862 425786 711098
rect 426022 710862 461786 711098
rect 462022 710862 497786 711098
rect 498022 710862 533786 711098
rect 534022 710862 569786 711098
rect 570022 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 29604 710838 30204 710840
rect 65604 710838 66204 710840
rect 101604 710838 102204 710840
rect 137604 710838 138204 710840
rect 173604 710838 174204 710840
rect 209604 710838 210204 710840
rect 245604 710838 246204 710840
rect 281604 710838 282204 710840
rect 317604 710838 318204 710840
rect 353604 710838 354204 710840
rect 389604 710838 390204 710840
rect 425604 710838 426204 710840
rect 461604 710838 462204 710840
rect 497604 710838 498204 710840
rect 533604 710838 534204 710840
rect 569604 710838 570204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 11604 710500 12204 710502
rect 47604 710500 48204 710502
rect 83604 710500 84204 710502
rect 119604 710500 120204 710502
rect 155604 710500 156204 710502
rect 191604 710500 192204 710502
rect 227604 710500 228204 710502
rect 263604 710500 264204 710502
rect 299604 710500 300204 710502
rect 335604 710500 336204 710502
rect 371604 710500 372204 710502
rect 407604 710500 408204 710502
rect 443604 710500 444204 710502
rect 479604 710500 480204 710502
rect 515604 710500 516204 710502
rect 551604 710500 552204 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 11786 710478
rect 12022 710242 47786 710478
rect 48022 710242 83786 710478
rect 84022 710242 119786 710478
rect 120022 710242 155786 710478
rect 156022 710242 191786 710478
rect 192022 710242 227786 710478
rect 228022 710242 263786 710478
rect 264022 710242 299786 710478
rect 300022 710242 335786 710478
rect 336022 710242 371786 710478
rect 372022 710242 407786 710478
rect 408022 710242 443786 710478
rect 444022 710242 479786 710478
rect 480022 710242 515786 710478
rect 516022 710242 551786 710478
rect 552022 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 11786 710158
rect 12022 709922 47786 710158
rect 48022 709922 83786 710158
rect 84022 709922 119786 710158
rect 120022 709922 155786 710158
rect 156022 709922 191786 710158
rect 192022 709922 227786 710158
rect 228022 709922 263786 710158
rect 264022 709922 299786 710158
rect 300022 709922 335786 710158
rect 336022 709922 371786 710158
rect 372022 709922 407786 710158
rect 408022 709922 443786 710158
rect 444022 709922 479786 710158
rect 480022 709922 515786 710158
rect 516022 709922 551786 710158
rect 552022 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 11604 709898 12204 709900
rect 47604 709898 48204 709900
rect 83604 709898 84204 709900
rect 119604 709898 120204 709900
rect 155604 709898 156204 709900
rect 191604 709898 192204 709900
rect 227604 709898 228204 709900
rect 263604 709898 264204 709900
rect 299604 709898 300204 709900
rect 335604 709898 336204 709900
rect 371604 709898 372204 709900
rect 407604 709898 408204 709900
rect 443604 709898 444204 709900
rect 479604 709898 480204 709900
rect 515604 709898 516204 709900
rect 551604 709898 552204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 26004 709560 26604 709562
rect 62004 709560 62604 709562
rect 98004 709560 98604 709562
rect 134004 709560 134604 709562
rect 170004 709560 170604 709562
rect 206004 709560 206604 709562
rect 242004 709560 242604 709562
rect 278004 709560 278604 709562
rect 314004 709560 314604 709562
rect 350004 709560 350604 709562
rect 386004 709560 386604 709562
rect 422004 709560 422604 709562
rect 458004 709560 458604 709562
rect 494004 709560 494604 709562
rect 530004 709560 530604 709562
rect 566004 709560 566604 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 26186 709538
rect 26422 709302 62186 709538
rect 62422 709302 98186 709538
rect 98422 709302 134186 709538
rect 134422 709302 170186 709538
rect 170422 709302 206186 709538
rect 206422 709302 242186 709538
rect 242422 709302 278186 709538
rect 278422 709302 314186 709538
rect 314422 709302 350186 709538
rect 350422 709302 386186 709538
rect 386422 709302 422186 709538
rect 422422 709302 458186 709538
rect 458422 709302 494186 709538
rect 494422 709302 530186 709538
rect 530422 709302 566186 709538
rect 566422 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 26186 709218
rect 26422 708982 62186 709218
rect 62422 708982 98186 709218
rect 98422 708982 134186 709218
rect 134422 708982 170186 709218
rect 170422 708982 206186 709218
rect 206422 708982 242186 709218
rect 242422 708982 278186 709218
rect 278422 708982 314186 709218
rect 314422 708982 350186 709218
rect 350422 708982 386186 709218
rect 386422 708982 422186 709218
rect 422422 708982 458186 709218
rect 458422 708982 494186 709218
rect 494422 708982 530186 709218
rect 530422 708982 566186 709218
rect 566422 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 26004 708958 26604 708960
rect 62004 708958 62604 708960
rect 98004 708958 98604 708960
rect 134004 708958 134604 708960
rect 170004 708958 170604 708960
rect 206004 708958 206604 708960
rect 242004 708958 242604 708960
rect 278004 708958 278604 708960
rect 314004 708958 314604 708960
rect 350004 708958 350604 708960
rect 386004 708958 386604 708960
rect 422004 708958 422604 708960
rect 458004 708958 458604 708960
rect 494004 708958 494604 708960
rect 530004 708958 530604 708960
rect 566004 708958 566604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 8004 708620 8604 708622
rect 44004 708620 44604 708622
rect 80004 708620 80604 708622
rect 116004 708620 116604 708622
rect 152004 708620 152604 708622
rect 188004 708620 188604 708622
rect 224004 708620 224604 708622
rect 260004 708620 260604 708622
rect 296004 708620 296604 708622
rect 332004 708620 332604 708622
rect 368004 708620 368604 708622
rect 404004 708620 404604 708622
rect 440004 708620 440604 708622
rect 476004 708620 476604 708622
rect 512004 708620 512604 708622
rect 548004 708620 548604 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 8186 708598
rect 8422 708362 44186 708598
rect 44422 708362 80186 708598
rect 80422 708362 116186 708598
rect 116422 708362 152186 708598
rect 152422 708362 188186 708598
rect 188422 708362 224186 708598
rect 224422 708362 260186 708598
rect 260422 708362 296186 708598
rect 296422 708362 332186 708598
rect 332422 708362 368186 708598
rect 368422 708362 404186 708598
rect 404422 708362 440186 708598
rect 440422 708362 476186 708598
rect 476422 708362 512186 708598
rect 512422 708362 548186 708598
rect 548422 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 8186 708278
rect 8422 708042 44186 708278
rect 44422 708042 80186 708278
rect 80422 708042 116186 708278
rect 116422 708042 152186 708278
rect 152422 708042 188186 708278
rect 188422 708042 224186 708278
rect 224422 708042 260186 708278
rect 260422 708042 296186 708278
rect 296422 708042 332186 708278
rect 332422 708042 368186 708278
rect 368422 708042 404186 708278
rect 404422 708042 440186 708278
rect 440422 708042 476186 708278
rect 476422 708042 512186 708278
rect 512422 708042 548186 708278
rect 548422 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 8004 708018 8604 708020
rect 44004 708018 44604 708020
rect 80004 708018 80604 708020
rect 116004 708018 116604 708020
rect 152004 708018 152604 708020
rect 188004 708018 188604 708020
rect 224004 708018 224604 708020
rect 260004 708018 260604 708020
rect 296004 708018 296604 708020
rect 332004 708018 332604 708020
rect 368004 708018 368604 708020
rect 404004 708018 404604 708020
rect 440004 708018 440604 708020
rect 476004 708018 476604 708020
rect 512004 708018 512604 708020
rect 548004 708018 548604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 22404 707680 23004 707682
rect 58404 707680 59004 707682
rect 94404 707680 95004 707682
rect 130404 707680 131004 707682
rect 166404 707680 167004 707682
rect 202404 707680 203004 707682
rect 238404 707680 239004 707682
rect 274404 707680 275004 707682
rect 310404 707680 311004 707682
rect 346404 707680 347004 707682
rect 382404 707680 383004 707682
rect 418404 707680 419004 707682
rect 454404 707680 455004 707682
rect 490404 707680 491004 707682
rect 526404 707680 527004 707682
rect 562404 707680 563004 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 22586 707658
rect 22822 707422 58586 707658
rect 58822 707422 94586 707658
rect 94822 707422 130586 707658
rect 130822 707422 166586 707658
rect 166822 707422 202586 707658
rect 202822 707422 238586 707658
rect 238822 707422 274586 707658
rect 274822 707422 310586 707658
rect 310822 707422 346586 707658
rect 346822 707422 382586 707658
rect 382822 707422 418586 707658
rect 418822 707422 454586 707658
rect 454822 707422 490586 707658
rect 490822 707422 526586 707658
rect 526822 707422 562586 707658
rect 562822 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 22586 707338
rect 22822 707102 58586 707338
rect 58822 707102 94586 707338
rect 94822 707102 130586 707338
rect 130822 707102 166586 707338
rect 166822 707102 202586 707338
rect 202822 707102 238586 707338
rect 238822 707102 274586 707338
rect 274822 707102 310586 707338
rect 310822 707102 346586 707338
rect 346822 707102 382586 707338
rect 382822 707102 418586 707338
rect 418822 707102 454586 707338
rect 454822 707102 490586 707338
rect 490822 707102 526586 707338
rect 526822 707102 562586 707338
rect 562822 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 22404 707078 23004 707080
rect 58404 707078 59004 707080
rect 94404 707078 95004 707080
rect 130404 707078 131004 707080
rect 166404 707078 167004 707080
rect 202404 707078 203004 707080
rect 238404 707078 239004 707080
rect 274404 707078 275004 707080
rect 310404 707078 311004 707080
rect 346404 707078 347004 707080
rect 382404 707078 383004 707080
rect 418404 707078 419004 707080
rect 454404 707078 455004 707080
rect 490404 707078 491004 707080
rect 526404 707078 527004 707080
rect 562404 707078 563004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 4404 706740 5004 706742
rect 40404 706740 41004 706742
rect 76404 706740 77004 706742
rect 112404 706740 113004 706742
rect 148404 706740 149004 706742
rect 184404 706740 185004 706742
rect 220404 706740 221004 706742
rect 256404 706740 257004 706742
rect 292404 706740 293004 706742
rect 328404 706740 329004 706742
rect 364404 706740 365004 706742
rect 400404 706740 401004 706742
rect 436404 706740 437004 706742
rect 472404 706740 473004 706742
rect 508404 706740 509004 706742
rect 544404 706740 545004 706742
rect 580404 706740 581004 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 4586 706718
rect 4822 706482 40586 706718
rect 40822 706482 76586 706718
rect 76822 706482 112586 706718
rect 112822 706482 148586 706718
rect 148822 706482 184586 706718
rect 184822 706482 220586 706718
rect 220822 706482 256586 706718
rect 256822 706482 292586 706718
rect 292822 706482 328586 706718
rect 328822 706482 364586 706718
rect 364822 706482 400586 706718
rect 400822 706482 436586 706718
rect 436822 706482 472586 706718
rect 472822 706482 508586 706718
rect 508822 706482 544586 706718
rect 544822 706482 580586 706718
rect 580822 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 4586 706398
rect 4822 706162 40586 706398
rect 40822 706162 76586 706398
rect 76822 706162 112586 706398
rect 112822 706162 148586 706398
rect 148822 706162 184586 706398
rect 184822 706162 220586 706398
rect 220822 706162 256586 706398
rect 256822 706162 292586 706398
rect 292822 706162 328586 706398
rect 328822 706162 364586 706398
rect 364822 706162 400586 706398
rect 400822 706162 436586 706398
rect 436822 706162 472586 706398
rect 472822 706162 508586 706398
rect 508822 706162 544586 706398
rect 544822 706162 580586 706398
rect 580822 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 4404 706138 5004 706140
rect 40404 706138 41004 706140
rect 76404 706138 77004 706140
rect 112404 706138 113004 706140
rect 148404 706138 149004 706140
rect 184404 706138 185004 706140
rect 220404 706138 221004 706140
rect 256404 706138 257004 706140
rect 292404 706138 293004 706140
rect 328404 706138 329004 706140
rect 364404 706138 365004 706140
rect 400404 706138 401004 706140
rect 436404 706138 437004 706140
rect 472404 706138 473004 706140
rect 508404 706138 509004 706140
rect 544404 706138 545004 706140
rect 580404 706138 581004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7636 697276 -7036 697278
rect 590960 697276 591560 697278
rect -8576 697254 480 697276
rect -8576 697018 -7454 697254
rect -7218 697018 480 697254
rect -8576 696934 480 697018
rect -8576 696698 -7454 696934
rect -7218 696698 480 696934
rect -8576 696676 480 696698
rect 583520 697254 592500 697276
rect 583520 697018 591142 697254
rect 591378 697018 592500 697254
rect 583520 696934 592500 697018
rect 583520 696698 591142 696934
rect 591378 696698 592500 696934
rect 583520 696676 592500 696698
rect -7636 696674 -7036 696676
rect 590960 696674 591560 696676
rect -5756 693676 -5156 693678
rect 589080 693676 589680 693678
rect -6696 693654 480 693676
rect -6696 693418 -5574 693654
rect -5338 693418 480 693654
rect -6696 693334 480 693418
rect -6696 693098 -5574 693334
rect -5338 693098 480 693334
rect -6696 693076 480 693098
rect 583520 693654 590620 693676
rect 583520 693418 589262 693654
rect 589498 693418 590620 693654
rect 583520 693334 590620 693418
rect 583520 693098 589262 693334
rect 589498 693098 590620 693334
rect 583520 693076 590620 693098
rect -5756 693074 -5156 693076
rect 589080 693074 589680 693076
rect -3876 690076 -3276 690078
rect 587200 690076 587800 690078
rect -4816 690054 480 690076
rect -4816 689818 -3694 690054
rect -3458 689818 480 690054
rect -4816 689734 480 689818
rect -4816 689498 -3694 689734
rect -3458 689498 480 689734
rect -4816 689476 480 689498
rect 583520 690054 588740 690076
rect 583520 689818 587382 690054
rect 587618 689818 588740 690054
rect 583520 689734 588740 689818
rect 583520 689498 587382 689734
rect 587618 689498 588740 689734
rect 583520 689476 588740 689498
rect -3876 689474 -3276 689476
rect 587200 689474 587800 689476
rect -1996 686476 -1396 686478
rect 585320 686476 585920 686478
rect -2936 686454 480 686476
rect -2936 686218 -1814 686454
rect -1578 686218 480 686454
rect -2936 686134 480 686218
rect -2936 685898 -1814 686134
rect -1578 685898 480 686134
rect -2936 685876 480 685898
rect 583520 686454 586860 686476
rect 583520 686218 585502 686454
rect 585738 686218 586860 686454
rect 583520 686134 586860 686218
rect 583520 685898 585502 686134
rect 585738 685898 586860 686134
rect 583520 685876 586860 685898
rect -1996 685874 -1396 685876
rect 585320 685874 585920 685876
rect -8576 679276 -7976 679278
rect 591900 679276 592500 679278
rect -8576 679254 480 679276
rect -8576 679018 -8394 679254
rect -8158 679018 480 679254
rect -8576 678934 480 679018
rect -8576 678698 -8394 678934
rect -8158 678698 480 678934
rect -8576 678676 480 678698
rect 583520 679254 592500 679276
rect 583520 679018 592082 679254
rect 592318 679018 592500 679254
rect 583520 678934 592500 679018
rect 583520 678698 592082 678934
rect 592318 678698 592500 678934
rect 583520 678676 592500 678698
rect -8576 678674 -7976 678676
rect 591900 678674 592500 678676
rect -6696 675676 -6096 675678
rect 590020 675676 590620 675678
rect -6696 675654 480 675676
rect -6696 675418 -6514 675654
rect -6278 675418 480 675654
rect -6696 675334 480 675418
rect -6696 675098 -6514 675334
rect -6278 675098 480 675334
rect -6696 675076 480 675098
rect 583520 675654 590620 675676
rect 583520 675418 590202 675654
rect 590438 675418 590620 675654
rect 583520 675334 590620 675418
rect 583520 675098 590202 675334
rect 590438 675098 590620 675334
rect 583520 675076 590620 675098
rect -6696 675074 -6096 675076
rect 590020 675074 590620 675076
rect -4816 672076 -4216 672078
rect 588140 672076 588740 672078
rect -4816 672054 480 672076
rect -4816 671818 -4634 672054
rect -4398 671818 480 672054
rect -4816 671734 480 671818
rect -4816 671498 -4634 671734
rect -4398 671498 480 671734
rect -4816 671476 480 671498
rect 583520 672054 588740 672076
rect 583520 671818 588322 672054
rect 588558 671818 588740 672054
rect 583520 671734 588740 671818
rect 583520 671498 588322 671734
rect 588558 671498 588740 671734
rect 583520 671476 588740 671498
rect -4816 671474 -4216 671476
rect 588140 671474 588740 671476
rect -2936 668476 -2336 668478
rect 586260 668476 586860 668478
rect -2936 668454 480 668476
rect -2936 668218 -2754 668454
rect -2518 668218 480 668454
rect -2936 668134 480 668218
rect -2936 667898 -2754 668134
rect -2518 667898 480 668134
rect -2936 667876 480 667898
rect 583520 668454 586860 668476
rect 583520 668218 586442 668454
rect 586678 668218 586860 668454
rect 583520 668134 586860 668218
rect 583520 667898 586442 668134
rect 586678 667898 586860 668134
rect 583520 667876 586860 667898
rect -2936 667874 -2336 667876
rect 586260 667874 586860 667876
rect -7636 661276 -7036 661278
rect 590960 661276 591560 661278
rect -8576 661254 480 661276
rect -8576 661018 -7454 661254
rect -7218 661018 480 661254
rect -8576 660934 480 661018
rect -8576 660698 -7454 660934
rect -7218 660698 480 660934
rect -8576 660676 480 660698
rect 583520 661254 592500 661276
rect 583520 661018 591142 661254
rect 591378 661018 592500 661254
rect 583520 660934 592500 661018
rect 583520 660698 591142 660934
rect 591378 660698 592500 660934
rect 583520 660676 592500 660698
rect -7636 660674 -7036 660676
rect 590960 660674 591560 660676
rect -5756 657676 -5156 657678
rect 589080 657676 589680 657678
rect -6696 657654 480 657676
rect -6696 657418 -5574 657654
rect -5338 657418 480 657654
rect -6696 657334 480 657418
rect -6696 657098 -5574 657334
rect -5338 657098 480 657334
rect -6696 657076 480 657098
rect 583520 657654 590620 657676
rect 583520 657418 589262 657654
rect 589498 657418 590620 657654
rect 583520 657334 590620 657418
rect 583520 657098 589262 657334
rect 589498 657098 590620 657334
rect 583520 657076 590620 657098
rect -5756 657074 -5156 657076
rect 589080 657074 589680 657076
rect -3876 654076 -3276 654078
rect 587200 654076 587800 654078
rect -4816 654054 480 654076
rect -4816 653818 -3694 654054
rect -3458 653818 480 654054
rect -4816 653734 480 653818
rect -4816 653498 -3694 653734
rect -3458 653498 480 653734
rect -4816 653476 480 653498
rect 583520 654054 588740 654076
rect 583520 653818 587382 654054
rect 587618 653818 588740 654054
rect 583520 653734 588740 653818
rect 583520 653498 587382 653734
rect 587618 653498 588740 653734
rect 583520 653476 588740 653498
rect -3876 653474 -3276 653476
rect 587200 653474 587800 653476
rect -1996 650476 -1396 650478
rect 585320 650476 585920 650478
rect -2936 650454 480 650476
rect -2936 650218 -1814 650454
rect -1578 650218 480 650454
rect -2936 650134 480 650218
rect -2936 649898 -1814 650134
rect -1578 649898 480 650134
rect -2936 649876 480 649898
rect 583520 650454 586860 650476
rect 583520 650218 585502 650454
rect 585738 650218 586860 650454
rect 583520 650134 586860 650218
rect 583520 649898 585502 650134
rect 585738 649898 586860 650134
rect 583520 649876 586860 649898
rect -1996 649874 -1396 649876
rect 585320 649874 585920 649876
rect -8576 643276 -7976 643278
rect 591900 643276 592500 643278
rect -8576 643254 480 643276
rect -8576 643018 -8394 643254
rect -8158 643018 480 643254
rect -8576 642934 480 643018
rect -8576 642698 -8394 642934
rect -8158 642698 480 642934
rect -8576 642676 480 642698
rect 583520 643254 592500 643276
rect 583520 643018 592082 643254
rect 592318 643018 592500 643254
rect 583520 642934 592500 643018
rect 583520 642698 592082 642934
rect 592318 642698 592500 642934
rect 583520 642676 592500 642698
rect -8576 642674 -7976 642676
rect 591900 642674 592500 642676
rect -6696 639676 -6096 639678
rect 590020 639676 590620 639678
rect -6696 639654 480 639676
rect -6696 639418 -6514 639654
rect -6278 639418 480 639654
rect -6696 639334 480 639418
rect -6696 639098 -6514 639334
rect -6278 639098 480 639334
rect -6696 639076 480 639098
rect 583520 639654 590620 639676
rect 583520 639418 590202 639654
rect 590438 639418 590620 639654
rect 583520 639334 590620 639418
rect 583520 639098 590202 639334
rect 590438 639098 590620 639334
rect 583520 639076 590620 639098
rect -6696 639074 -6096 639076
rect 590020 639074 590620 639076
rect -4816 636076 -4216 636078
rect 588140 636076 588740 636078
rect -4816 636054 480 636076
rect -4816 635818 -4634 636054
rect -4398 635818 480 636054
rect -4816 635734 480 635818
rect -4816 635498 -4634 635734
rect -4398 635498 480 635734
rect -4816 635476 480 635498
rect 583520 636054 588740 636076
rect 583520 635818 588322 636054
rect 588558 635818 588740 636054
rect 583520 635734 588740 635818
rect 583520 635498 588322 635734
rect 588558 635498 588740 635734
rect 583520 635476 588740 635498
rect -4816 635474 -4216 635476
rect 588140 635474 588740 635476
rect -2936 632476 -2336 632478
rect 586260 632476 586860 632478
rect -2936 632454 480 632476
rect -2936 632218 -2754 632454
rect -2518 632218 480 632454
rect -2936 632134 480 632218
rect -2936 631898 -2754 632134
rect -2518 631898 480 632134
rect -2936 631876 480 631898
rect 545212 632454 586860 632476
rect 545212 632450 586442 632454
rect 545212 632214 545562 632450
rect 545798 632218 586442 632450
rect 586678 632218 586860 632454
rect 545798 632214 586860 632218
rect 545212 632134 586860 632214
rect 545212 632130 586442 632134
rect 545212 631894 545562 632130
rect 545798 631898 586442 632130
rect 586678 631898 586860 632134
rect 545798 631894 586860 631898
rect 545212 631876 586860 631894
rect -2936 631874 -2336 631876
rect 545224 631868 546170 631876
rect 586260 631874 586860 631876
rect -7636 625276 -7036 625278
rect 590960 625276 591560 625278
rect -8576 625254 480 625276
rect -8576 625018 -7454 625254
rect -7218 625018 480 625254
rect -8576 624934 480 625018
rect -8576 624698 -7454 624934
rect -7218 624698 480 624934
rect -8576 624676 480 624698
rect 583520 625254 592500 625276
rect 583520 625018 591142 625254
rect 591378 625018 592500 625254
rect 583520 624934 592500 625018
rect 583520 624698 591142 624934
rect 591378 624698 592500 624934
rect 583520 624676 592500 624698
rect -7636 624674 -7036 624676
rect 590960 624674 591560 624676
rect -5756 621676 -5156 621678
rect 589080 621676 589680 621678
rect -6696 621654 480 621676
rect -6696 621418 -5574 621654
rect -5338 621418 480 621654
rect -6696 621334 480 621418
rect -6696 621098 -5574 621334
rect -5338 621098 480 621334
rect -6696 621076 480 621098
rect 583520 621654 590620 621676
rect 583520 621418 589262 621654
rect 589498 621418 590620 621654
rect 583520 621334 590620 621418
rect 583520 621098 589262 621334
rect 589498 621098 590620 621334
rect 583520 621076 590620 621098
rect -5756 621074 -5156 621076
rect 589080 621074 589680 621076
rect -3876 618076 -3276 618078
rect 587200 618076 587800 618078
rect -4816 618054 480 618076
rect -4816 617818 -3694 618054
rect -3458 617818 480 618054
rect -4816 617734 480 617818
rect -4816 617498 -3694 617734
rect -3458 617498 480 617734
rect -4816 617476 480 617498
rect 583520 618054 588740 618076
rect 583520 617818 587382 618054
rect 587618 617818 588740 618054
rect 583520 617734 588740 617818
rect 583520 617498 587382 617734
rect 587618 617498 588740 617734
rect 583520 617476 588740 617498
rect -3876 617474 -3276 617476
rect 587200 617474 587800 617476
rect -1996 614476 -1396 614478
rect 585320 614476 585920 614478
rect -2936 614454 480 614476
rect -2936 614218 -1814 614454
rect -1578 614218 480 614454
rect -2936 614134 480 614218
rect -2936 613898 -1814 614134
rect -1578 613898 480 614134
rect -2936 613876 480 613898
rect 583508 614454 586860 614476
rect 583508 614218 585502 614454
rect 585738 614218 586860 614454
rect 583508 614134 586860 614218
rect 583508 613898 585502 614134
rect 585738 613898 586860 614134
rect 583508 613876 586860 613898
rect -1996 613874 -1396 613876
rect 585320 613874 585920 613876
rect -8576 607276 -7976 607278
rect 591900 607276 592500 607278
rect -8576 607254 480 607276
rect -8576 607018 -8394 607254
rect -8158 607018 480 607254
rect -8576 606934 480 607018
rect -8576 606698 -8394 606934
rect -8158 606698 480 606934
rect -8576 606676 480 606698
rect 583520 607254 592500 607276
rect 583520 607018 592082 607254
rect 592318 607018 592500 607254
rect 583520 606934 592500 607018
rect 583520 606698 592082 606934
rect 592318 606698 592500 606934
rect 583520 606676 592500 606698
rect -8576 606674 -7976 606676
rect 591900 606674 592500 606676
rect -6696 603676 -6096 603678
rect 590020 603676 590620 603678
rect -6696 603654 480 603676
rect -6696 603418 -6514 603654
rect -6278 603418 480 603654
rect -6696 603334 480 603418
rect -6696 603098 -6514 603334
rect -6278 603098 480 603334
rect -6696 603076 480 603098
rect 583520 603654 590620 603676
rect 583520 603418 590202 603654
rect 590438 603418 590620 603654
rect 583520 603334 590620 603418
rect 583520 603098 590202 603334
rect 590438 603098 590620 603334
rect 583520 603076 590620 603098
rect -6696 603074 -6096 603076
rect 590020 603074 590620 603076
rect -4816 600076 -4216 600078
rect 588140 600076 588740 600078
rect -4816 600054 480 600076
rect -4816 599818 -4634 600054
rect -4398 599818 480 600054
rect -4816 599734 480 599818
rect -4816 599498 -4634 599734
rect -4398 599498 480 599734
rect -4816 599476 480 599498
rect 583520 600054 588740 600076
rect 583520 599818 588322 600054
rect 588558 599818 588740 600054
rect 583520 599734 588740 599818
rect 583520 599498 588322 599734
rect 588558 599498 588740 599734
rect 583520 599476 588740 599498
rect -4816 599474 -4216 599476
rect 588140 599474 588740 599476
rect -2936 596476 -2336 596478
rect 35324 596476 35924 596478
rect 586260 596476 586860 596478
rect -2936 596474 36014 596476
rect -2936 596454 36016 596474
rect -2936 596218 -2754 596454
rect -2518 596218 35506 596454
rect 35742 596218 36016 596454
rect -2936 596134 36016 596218
rect -2936 595898 -2754 596134
rect -2518 595898 35506 596134
rect 35742 595898 36016 596134
rect -2936 595876 36016 595898
rect 583520 596454 586860 596476
rect 583520 596218 586442 596454
rect 586678 596218 586860 596454
rect 583520 596134 586860 596218
rect 583520 595898 586442 596134
rect 586678 595898 586860 596134
rect 583520 595876 586860 595898
rect -2936 595874 -2336 595876
rect 35254 595874 36016 595876
rect 586260 595874 586860 595876
rect -7636 589276 -7036 589278
rect 590960 589276 591560 589278
rect -8576 589254 480 589276
rect -8576 589018 -7454 589254
rect -7218 589018 480 589254
rect -8576 588934 480 589018
rect -8576 588698 -7454 588934
rect -7218 588698 480 588934
rect -8576 588676 480 588698
rect 583520 589254 592500 589276
rect 583520 589018 591142 589254
rect 591378 589018 592500 589254
rect 583520 588934 592500 589018
rect 583520 588698 591142 588934
rect 591378 588698 592500 588934
rect 583520 588676 592500 588698
rect -7636 588674 -7036 588676
rect 590960 588674 591560 588676
rect -5756 585676 -5156 585678
rect 589080 585676 589680 585678
rect -6696 585654 480 585676
rect -6696 585418 -5574 585654
rect -5338 585418 480 585654
rect -6696 585334 480 585418
rect -6696 585098 -5574 585334
rect -5338 585098 480 585334
rect -6696 585076 480 585098
rect 583520 585654 590620 585676
rect 583520 585418 589262 585654
rect 589498 585418 590620 585654
rect 583520 585334 590620 585418
rect 583520 585098 589262 585334
rect 589498 585098 590620 585334
rect 583520 585076 590620 585098
rect -5756 585074 -5156 585076
rect 589080 585074 589680 585076
rect -3876 582076 -3276 582078
rect 587200 582076 587800 582078
rect -4816 582054 480 582076
rect -4816 581818 -3694 582054
rect -3458 581818 480 582054
rect -4816 581734 480 581818
rect -4816 581498 -3694 581734
rect -3458 581498 480 581734
rect -4816 581476 480 581498
rect 583520 582054 588740 582076
rect 583520 581818 587382 582054
rect 587618 581818 588740 582054
rect 583520 581734 588740 581818
rect 583520 581498 587382 581734
rect 587618 581498 588740 581734
rect 583520 581476 588740 581498
rect -3876 581474 -3276 581476
rect 587200 581474 587800 581476
rect -1996 578476 -1396 578478
rect 585320 578476 585920 578478
rect -2936 578454 480 578476
rect -2936 578218 -1814 578454
rect -1578 578218 480 578454
rect -2936 578134 480 578218
rect -2936 577898 -1814 578134
rect -1578 577898 480 578134
rect -2936 577876 480 577898
rect 545616 578454 586860 578476
rect 545616 578452 585502 578454
rect 545616 578216 545990 578452
rect 546226 578218 585502 578452
rect 585738 578218 586860 578454
rect 546226 578216 586860 578218
rect 545616 578134 586860 578216
rect 545616 578132 585502 578134
rect 545616 577896 545990 578132
rect 546226 577898 585502 578132
rect 585738 577898 586860 578134
rect 546226 577896 586860 577898
rect 545616 577876 586860 577896
rect -1996 577874 -1396 577876
rect 545738 577872 546642 577876
rect 585320 577874 585920 577876
rect -8576 571276 -7976 571278
rect 591900 571276 592500 571278
rect -8576 571254 480 571276
rect -8576 571018 -8394 571254
rect -8158 571018 480 571254
rect -8576 570934 480 571018
rect -8576 570698 -8394 570934
rect -8158 570698 480 570934
rect -8576 570676 480 570698
rect 583520 571254 592500 571276
rect 583520 571018 592082 571254
rect 592318 571018 592500 571254
rect 583520 570934 592500 571018
rect 583520 570698 592082 570934
rect 592318 570698 592500 570934
rect 583520 570676 592500 570698
rect -8576 570674 -7976 570676
rect 591900 570674 592500 570676
rect -6696 567676 -6096 567678
rect 590020 567676 590620 567678
rect -6696 567654 480 567676
rect -6696 567418 -6514 567654
rect -6278 567418 480 567654
rect -6696 567334 480 567418
rect -6696 567098 -6514 567334
rect -6278 567098 480 567334
rect -6696 567076 480 567098
rect 583520 567654 590620 567676
rect 583520 567418 590202 567654
rect 590438 567418 590620 567654
rect 583520 567334 590620 567418
rect 583520 567098 590202 567334
rect 590438 567098 590620 567334
rect 583520 567076 590620 567098
rect -6696 567074 -6096 567076
rect 590020 567074 590620 567076
rect -4816 564076 -4216 564078
rect 588140 564076 588740 564078
rect -4816 564054 480 564076
rect -4816 563818 -4634 564054
rect -4398 563818 480 564054
rect -4816 563734 480 563818
rect -4816 563498 -4634 563734
rect -4398 563498 480 563734
rect -4816 563476 480 563498
rect 583520 564054 588740 564076
rect 583520 563818 588322 564054
rect 588558 563818 588740 564054
rect 583520 563734 588740 563818
rect 583520 563498 588322 563734
rect 588558 563498 588740 563734
rect 583520 563476 588740 563498
rect -4816 563474 -4216 563476
rect 588140 563474 588740 563476
rect -2936 560476 -2336 560478
rect 586260 560476 586860 560478
rect -2936 560454 480 560476
rect -2936 560218 -2754 560454
rect -2518 560218 480 560454
rect -2936 560134 480 560218
rect -2936 559898 -2754 560134
rect -2518 559898 480 560134
rect -2936 559876 480 559898
rect 583512 560454 586860 560476
rect 583512 560218 586442 560454
rect 586678 560218 586860 560454
rect 583512 560134 586860 560218
rect 583512 559898 586442 560134
rect 586678 559898 586860 560134
rect 583512 559876 586860 559898
rect -2936 559874 -2336 559876
rect 586260 559874 586860 559876
rect -7636 553276 -7036 553278
rect 590960 553276 591560 553278
rect -8576 553254 480 553276
rect -8576 553018 -7454 553254
rect -7218 553018 480 553254
rect -8576 552934 480 553018
rect -8576 552698 -7454 552934
rect -7218 552698 480 552934
rect -8576 552676 480 552698
rect 583520 553254 592500 553276
rect 583520 553018 591142 553254
rect 591378 553018 592500 553254
rect 583520 552934 592500 553018
rect 583520 552698 591142 552934
rect 591378 552698 592500 552934
rect 583520 552676 592500 552698
rect -7636 552674 -7036 552676
rect 590960 552674 591560 552676
rect -5756 549676 -5156 549678
rect 589080 549676 589680 549678
rect -6696 549654 480 549676
rect -6696 549418 -5574 549654
rect -5338 549418 480 549654
rect -6696 549334 480 549418
rect -6696 549098 -5574 549334
rect -5338 549098 480 549334
rect -6696 549076 480 549098
rect 583520 549654 590620 549676
rect 583520 549418 589262 549654
rect 589498 549418 590620 549654
rect 583520 549334 590620 549418
rect 583520 549098 589262 549334
rect 589498 549098 590620 549334
rect 583520 549076 590620 549098
rect -5756 549074 -5156 549076
rect 589080 549074 589680 549076
rect -3876 546076 -3276 546078
rect 587200 546076 587800 546078
rect -4816 546054 480 546076
rect -4816 545818 -3694 546054
rect -3458 545818 480 546054
rect -4816 545734 480 545818
rect -4816 545498 -3694 545734
rect -3458 545498 480 545734
rect -4816 545476 480 545498
rect 583520 546054 588740 546076
rect 583520 545818 587382 546054
rect 587618 545818 588740 546054
rect 583520 545734 588740 545818
rect 583520 545498 587382 545734
rect 587618 545498 588740 545734
rect 583520 545476 588740 545498
rect -3876 545474 -3276 545476
rect 587200 545474 587800 545476
rect -1996 542476 -1396 542478
rect 585320 542476 585920 542478
rect -2936 542454 480 542476
rect -2936 542218 -1814 542454
rect -1578 542218 480 542454
rect -2936 542134 480 542218
rect -2936 541898 -1814 542134
rect -1578 541898 480 542134
rect -2936 541876 480 541898
rect 583520 542454 586860 542476
rect 583520 542218 585502 542454
rect 585738 542218 586860 542454
rect 583520 542134 586860 542218
rect 583520 541898 585502 542134
rect 585738 541898 586860 542134
rect 583520 541876 586860 541898
rect -1996 541874 -1396 541876
rect 585320 541874 585920 541876
rect -8576 535276 -7976 535278
rect 591900 535276 592500 535278
rect -8576 535254 480 535276
rect -8576 535018 -8394 535254
rect -8158 535018 480 535254
rect -8576 534934 480 535018
rect -8576 534698 -8394 534934
rect -8158 534698 480 534934
rect -8576 534676 480 534698
rect 583520 535254 592500 535276
rect 583520 535018 592082 535254
rect 592318 535018 592500 535254
rect 583520 534934 592500 535018
rect 583520 534698 592082 534934
rect 592318 534698 592500 534934
rect 583520 534676 592500 534698
rect -8576 534674 -7976 534676
rect 591900 534674 592500 534676
rect -6696 531676 -6096 531678
rect 590020 531676 590620 531678
rect -6696 531654 480 531676
rect -6696 531418 -6514 531654
rect -6278 531418 480 531654
rect -6696 531334 480 531418
rect -6696 531098 -6514 531334
rect -6278 531098 480 531334
rect -6696 531076 480 531098
rect 583520 531654 590620 531676
rect 583520 531418 590202 531654
rect 590438 531418 590620 531654
rect 583520 531334 590620 531418
rect 583520 531098 590202 531334
rect 590438 531098 590620 531334
rect 583520 531076 590620 531098
rect -6696 531074 -6096 531076
rect 590020 531074 590620 531076
rect -4816 528076 -4216 528078
rect 588140 528076 588740 528078
rect -4816 528054 480 528076
rect -4816 527818 -4634 528054
rect -4398 527818 480 528054
rect -4816 527734 480 527818
rect -4816 527498 -4634 527734
rect -4398 527498 480 527734
rect -4816 527476 480 527498
rect 583520 528054 588740 528076
rect 583520 527818 588322 528054
rect 588558 527818 588740 528054
rect 583520 527734 588740 527818
rect 583520 527498 588322 527734
rect 588558 527498 588740 527734
rect 583520 527476 588740 527498
rect -4816 527474 -4216 527476
rect 588140 527474 588740 527476
rect -2936 524476 -2336 524478
rect 586260 524476 586860 524478
rect -2936 524454 480 524476
rect -2936 524218 -2754 524454
rect -2518 524218 480 524454
rect -2936 524134 480 524218
rect -2936 523898 -2754 524134
rect -2518 523898 480 524134
rect -2936 523876 480 523898
rect 583520 524454 586860 524476
rect 583520 524218 586442 524454
rect 586678 524218 586860 524454
rect 583520 524134 586860 524218
rect 583520 523898 586442 524134
rect 586678 523898 586860 524134
rect 583520 523876 586860 523898
rect -2936 523874 -2336 523876
rect 586260 523874 586860 523876
rect -7636 517276 -7036 517278
rect 590960 517276 591560 517278
rect -8576 517254 480 517276
rect -8576 517018 -7454 517254
rect -7218 517018 480 517254
rect -8576 516934 480 517018
rect -8576 516698 -7454 516934
rect -7218 516698 480 516934
rect -8576 516676 480 516698
rect 583520 517254 592500 517276
rect 583520 517018 591142 517254
rect 591378 517018 592500 517254
rect 583520 516934 592500 517018
rect 583520 516698 591142 516934
rect 591378 516698 592500 516934
rect 583520 516676 592500 516698
rect -7636 516674 -7036 516676
rect 590960 516674 591560 516676
rect -5756 513676 -5156 513678
rect 589080 513676 589680 513678
rect -6696 513654 480 513676
rect -6696 513418 -5574 513654
rect -5338 513418 480 513654
rect -6696 513334 480 513418
rect -6696 513098 -5574 513334
rect -5338 513098 480 513334
rect -6696 513076 480 513098
rect 583520 513654 590620 513676
rect 583520 513418 589262 513654
rect 589498 513418 590620 513654
rect 583520 513334 590620 513418
rect 583520 513098 589262 513334
rect 589498 513098 590620 513334
rect 583520 513076 590620 513098
rect -5756 513074 -5156 513076
rect 589080 513074 589680 513076
rect -3876 510076 -3276 510078
rect 587200 510076 587800 510078
rect -4816 510054 480 510076
rect -4816 509818 -3694 510054
rect -3458 509818 480 510054
rect -4816 509734 480 509818
rect -4816 509498 -3694 509734
rect -3458 509498 480 509734
rect -4816 509476 480 509498
rect 583520 510054 588740 510076
rect 583520 509818 587382 510054
rect 587618 509818 588740 510054
rect 583520 509734 588740 509818
rect 583520 509498 587382 509734
rect 587618 509498 588740 509734
rect 583520 509476 588740 509498
rect -3876 509474 -3276 509476
rect 587200 509474 587800 509476
rect -1996 506476 -1396 506478
rect 585320 506476 585920 506478
rect -2936 506454 480 506476
rect -2936 506218 -1814 506454
rect -1578 506218 480 506454
rect -2936 506134 480 506218
rect -2936 505898 -1814 506134
rect -1578 505898 480 506134
rect -2936 505876 480 505898
rect 583520 506454 586860 506476
rect 583520 506218 585502 506454
rect 585738 506218 586860 506454
rect 583520 506134 586860 506218
rect 583520 505898 585502 506134
rect 585738 505898 586860 506134
rect 583520 505876 586860 505898
rect -1996 505874 -1396 505876
rect 585320 505874 585920 505876
rect -8576 499276 -7976 499278
rect 591900 499276 592500 499278
rect -8576 499254 480 499276
rect -8576 499018 -8394 499254
rect -8158 499018 480 499254
rect -8576 498934 480 499018
rect -8576 498698 -8394 498934
rect -8158 498698 480 498934
rect -8576 498676 480 498698
rect 583520 499254 592500 499276
rect 583520 499018 592082 499254
rect 592318 499018 592500 499254
rect 583520 498934 592500 499018
rect 583520 498698 592082 498934
rect 592318 498698 592500 498934
rect 583520 498676 592500 498698
rect -8576 498674 -7976 498676
rect 591900 498674 592500 498676
rect -6696 495676 -6096 495678
rect 590020 495676 590620 495678
rect -6696 495654 480 495676
rect -6696 495418 -6514 495654
rect -6278 495418 480 495654
rect -6696 495334 480 495418
rect -6696 495098 -6514 495334
rect -6278 495098 480 495334
rect -6696 495076 480 495098
rect 583520 495654 590620 495676
rect 583520 495418 590202 495654
rect 590438 495418 590620 495654
rect 583520 495334 590620 495418
rect 583520 495098 590202 495334
rect 590438 495098 590620 495334
rect 583520 495076 590620 495098
rect -6696 495074 -6096 495076
rect 590020 495074 590620 495076
rect -4816 492076 -4216 492078
rect 588140 492076 588740 492078
rect -4816 492054 480 492076
rect -4816 491818 -4634 492054
rect -4398 491818 480 492054
rect -4816 491734 480 491818
rect -4816 491498 -4634 491734
rect -4398 491498 480 491734
rect -4816 491476 480 491498
rect 583520 492054 588740 492076
rect 583520 491818 588322 492054
rect 588558 491818 588740 492054
rect 583520 491734 588740 491818
rect 583520 491498 588322 491734
rect 588558 491498 588740 491734
rect 583520 491476 588740 491498
rect -4816 491474 -4216 491476
rect 588140 491474 588740 491476
rect -2936 488476 -2336 488478
rect 586260 488476 586860 488478
rect -2936 488454 480 488476
rect -2936 488218 -2754 488454
rect -2518 488218 480 488454
rect -2936 488134 480 488218
rect -2936 487898 -2754 488134
rect -2518 487898 480 488134
rect -2936 487876 480 487898
rect 583520 488454 586860 488476
rect 583520 488218 586442 488454
rect 586678 488218 586860 488454
rect 583520 488134 586860 488218
rect 583520 487898 586442 488134
rect 586678 487898 586860 488134
rect 583520 487876 586860 487898
rect -2936 487874 -2336 487876
rect 586260 487874 586860 487876
rect -7636 481276 -7036 481278
rect 590960 481276 591560 481278
rect -8576 481254 480 481276
rect -8576 481018 -7454 481254
rect -7218 481018 480 481254
rect -8576 480934 480 481018
rect -8576 480698 -7454 480934
rect -7218 480698 480 480934
rect -8576 480676 480 480698
rect 583520 481254 592500 481276
rect 583520 481018 591142 481254
rect 591378 481018 592500 481254
rect 583520 480934 592500 481018
rect 583520 480698 591142 480934
rect 591378 480698 592500 480934
rect 583520 480676 592500 480698
rect -7636 480674 -7036 480676
rect 590960 480674 591560 480676
rect -5756 477676 -5156 477678
rect 589080 477676 589680 477678
rect -6696 477654 480 477676
rect -6696 477418 -5574 477654
rect -5338 477418 480 477654
rect -6696 477334 480 477418
rect -6696 477098 -5574 477334
rect -5338 477098 480 477334
rect -6696 477076 480 477098
rect 583520 477654 590620 477676
rect 583520 477418 589262 477654
rect 589498 477418 590620 477654
rect 583520 477334 590620 477418
rect 583520 477098 589262 477334
rect 589498 477098 590620 477334
rect 583520 477076 590620 477098
rect -5756 477074 -5156 477076
rect 589080 477074 589680 477076
rect -3876 474076 -3276 474078
rect 587200 474076 587800 474078
rect -4816 474054 480 474076
rect -4816 473818 -3694 474054
rect -3458 473818 480 474054
rect -4816 473734 480 473818
rect -4816 473498 -3694 473734
rect -3458 473498 480 473734
rect -4816 473476 480 473498
rect 583520 474054 588740 474076
rect 583520 473818 587382 474054
rect 587618 473818 588740 474054
rect 583520 473734 588740 473818
rect 583520 473498 587382 473734
rect 587618 473498 588740 473734
rect 583520 473476 588740 473498
rect -3876 473474 -3276 473476
rect 587200 473474 587800 473476
rect -1996 470476 -1396 470478
rect 34418 470476 35018 470478
rect 585320 470476 585920 470478
rect -2936 470454 35018 470476
rect -2936 470218 -1814 470454
rect -1578 470218 34600 470454
rect 34836 470218 35018 470454
rect -2936 470134 35018 470218
rect -2936 469898 -1814 470134
rect -1578 469898 34600 470134
rect 34836 469898 35018 470134
rect -2936 469876 35018 469898
rect 583520 470454 586860 470476
rect 583520 470218 585502 470454
rect 585738 470218 586860 470454
rect 583520 470134 586860 470218
rect 583520 469898 585502 470134
rect 585738 469898 586860 470134
rect 583520 469876 586860 469898
rect -1996 469874 -1396 469876
rect 34418 469874 35018 469876
rect 585320 469874 585920 469876
rect -8576 463276 -7976 463278
rect 591900 463276 592500 463278
rect -8576 463254 480 463276
rect -8576 463018 -8394 463254
rect -8158 463018 480 463254
rect -8576 462934 480 463018
rect -8576 462698 -8394 462934
rect -8158 462698 480 462934
rect -8576 462676 480 462698
rect 583520 463254 592500 463276
rect 583520 463018 592082 463254
rect 592318 463018 592500 463254
rect 583520 462934 592500 463018
rect 583520 462698 592082 462934
rect 592318 462698 592500 462934
rect 583520 462676 592500 462698
rect -8576 462674 -7976 462676
rect 591900 462674 592500 462676
rect -6696 459676 -6096 459678
rect 590020 459676 590620 459678
rect -6696 459654 480 459676
rect -6696 459418 -6514 459654
rect -6278 459418 480 459654
rect -6696 459334 480 459418
rect -6696 459098 -6514 459334
rect -6278 459098 480 459334
rect -6696 459076 480 459098
rect 583520 459654 590620 459676
rect 583520 459418 590202 459654
rect 590438 459418 590620 459654
rect 583520 459334 590620 459418
rect 583520 459098 590202 459334
rect 590438 459098 590620 459334
rect 583520 459076 590620 459098
rect -6696 459074 -6096 459076
rect 590020 459074 590620 459076
rect -4816 456076 -4216 456078
rect 588140 456076 588740 456078
rect -4816 456054 480 456076
rect -4816 455818 -4634 456054
rect -4398 455818 480 456054
rect -4816 455734 480 455818
rect -4816 455498 -4634 455734
rect -4398 455498 480 455734
rect -4816 455476 480 455498
rect 583520 456054 588740 456076
rect 583520 455818 588322 456054
rect 588558 455818 588740 456054
rect 583520 455734 588740 455818
rect 583520 455498 588322 455734
rect 588558 455498 588740 455734
rect 583520 455476 588740 455498
rect -4816 455474 -4216 455476
rect 588140 455474 588740 455476
rect -2936 452476 -2336 452478
rect 586260 452476 586860 452478
rect -2936 452454 480 452476
rect -2936 452218 -2754 452454
rect -2518 452218 480 452454
rect -2936 452134 480 452218
rect -2936 451898 -2754 452134
rect -2518 451898 480 452134
rect -2936 451876 480 451898
rect 583520 452454 586860 452476
rect 583520 452218 586442 452454
rect 586678 452218 586860 452454
rect 583520 452134 586860 452218
rect 583520 451898 586442 452134
rect 586678 451898 586860 452134
rect 583520 451876 586860 451898
rect -2936 451874 -2336 451876
rect 586260 451874 586860 451876
rect -7636 445276 -7036 445278
rect 590960 445276 591560 445278
rect -8576 445254 480 445276
rect -8576 445018 -7454 445254
rect -7218 445018 480 445254
rect -8576 444934 480 445018
rect -8576 444698 -7454 444934
rect -7218 444698 480 444934
rect -8576 444676 480 444698
rect 583520 445254 592500 445276
rect 583520 445018 591142 445254
rect 591378 445018 592500 445254
rect 583520 444934 592500 445018
rect 583520 444698 591142 444934
rect 591378 444698 592500 444934
rect 583520 444676 592500 444698
rect -7636 444674 -7036 444676
rect 590960 444674 591560 444676
rect -5756 441676 -5156 441678
rect 589080 441676 589680 441678
rect -6696 441654 480 441676
rect -6696 441418 -5574 441654
rect -5338 441418 480 441654
rect -6696 441334 480 441418
rect -6696 441098 -5574 441334
rect -5338 441098 480 441334
rect -6696 441076 480 441098
rect 583520 441654 590620 441676
rect 583520 441418 589262 441654
rect 589498 441418 590620 441654
rect 583520 441334 590620 441418
rect 583520 441098 589262 441334
rect 589498 441098 590620 441334
rect 583520 441076 590620 441098
rect -5756 441074 -5156 441076
rect 589080 441074 589680 441076
rect -3876 438076 -3276 438078
rect 587200 438076 587800 438078
rect -4816 438054 480 438076
rect -4816 437818 -3694 438054
rect -3458 437818 480 438054
rect -4816 437734 480 437818
rect -4816 437498 -3694 437734
rect -3458 437498 480 437734
rect -4816 437476 480 437498
rect 583520 438054 588740 438076
rect 583520 437818 587382 438054
rect 587618 437818 588740 438054
rect 583520 437734 588740 437818
rect 583520 437498 587382 437734
rect 587618 437498 588740 437734
rect 583520 437476 588740 437498
rect -3876 437474 -3276 437476
rect 587200 437474 587800 437476
rect -1996 434476 -1396 434478
rect 585320 434476 585920 434478
rect -2936 434454 480 434476
rect -2936 434218 -1814 434454
rect -1578 434218 480 434454
rect -2936 434134 480 434218
rect -2936 433898 -1814 434134
rect -1578 433898 480 434134
rect -2936 433876 480 433898
rect 583496 434454 586860 434476
rect 583496 434218 585502 434454
rect 585738 434218 586860 434454
rect 583496 434134 586860 434218
rect 583496 433898 585502 434134
rect 585738 433898 586860 434134
rect 583496 433876 586860 433898
rect -1996 433874 -1396 433876
rect 585320 433874 585920 433876
rect -8576 427276 -7976 427278
rect 591900 427276 592500 427278
rect -8576 427254 480 427276
rect -8576 427018 -8394 427254
rect -8158 427018 480 427254
rect -8576 426934 480 427018
rect -8576 426698 -8394 426934
rect -8158 426698 480 426934
rect -8576 426676 480 426698
rect 583520 427254 592500 427276
rect 583520 427018 592082 427254
rect 592318 427018 592500 427254
rect 583520 426934 592500 427018
rect 583520 426698 592082 426934
rect 592318 426698 592500 426934
rect 583520 426676 592500 426698
rect -8576 426674 -7976 426676
rect 591900 426674 592500 426676
rect -6696 423676 -6096 423678
rect 590020 423676 590620 423678
rect -6696 423654 480 423676
rect -6696 423418 -6514 423654
rect -6278 423418 480 423654
rect -6696 423334 480 423418
rect -6696 423098 -6514 423334
rect -6278 423098 480 423334
rect -6696 423076 480 423098
rect 583520 423654 590620 423676
rect 583520 423418 590202 423654
rect 590438 423418 590620 423654
rect 583520 423334 590620 423418
rect 583520 423098 590202 423334
rect 590438 423098 590620 423334
rect 583520 423076 590620 423098
rect -6696 423074 -6096 423076
rect 590020 423074 590620 423076
rect -4816 420076 -4216 420078
rect 588140 420076 588740 420078
rect -4816 420054 480 420076
rect -4816 419818 -4634 420054
rect -4398 419818 480 420054
rect -4816 419734 480 419818
rect -4816 419498 -4634 419734
rect -4398 419498 480 419734
rect -4816 419476 480 419498
rect 583520 420054 588740 420076
rect 583520 419818 588322 420054
rect 588558 419818 588740 420054
rect 583520 419734 588740 419818
rect 583520 419498 588322 419734
rect 588558 419498 588740 419734
rect 583520 419476 588740 419498
rect -4816 419474 -4216 419476
rect 588140 419474 588740 419476
rect 34852 416478 35452 416480
rect -2936 416476 -2336 416478
rect 34830 416476 35452 416478
rect 545260 416476 546216 416482
rect 586260 416476 586860 416478
rect -2936 416456 35610 416476
rect -2936 416454 35034 416456
rect -2936 416218 -2754 416454
rect -2518 416220 35034 416454
rect 35270 416220 35610 416456
rect -2518 416218 35610 416220
rect -2936 416136 35610 416218
rect -2936 416134 35034 416136
rect -2936 415898 -2754 416134
rect -2518 415900 35034 416134
rect 35270 415900 35610 416136
rect -2518 415898 35610 415900
rect -2936 415876 35610 415898
rect 545234 416454 586860 416476
rect 545234 416446 586442 416454
rect 545234 416210 545560 416446
rect 545796 416218 586442 416446
rect 586678 416218 586860 416454
rect 545796 416210 586860 416218
rect 545234 416134 586860 416210
rect 545234 416126 586442 416134
rect 545234 415890 545560 416126
rect 545796 415898 586442 416126
rect 586678 415898 586860 416134
rect 545796 415890 586860 415898
rect 545234 415876 586860 415890
rect -2936 415874 -2336 415876
rect 545260 415864 546116 415876
rect 586260 415874 586860 415876
rect -7636 409276 -7036 409278
rect 590960 409276 591560 409278
rect -8576 409254 480 409276
rect -8576 409018 -7454 409254
rect -7218 409018 480 409254
rect -8576 408934 480 409018
rect -8576 408698 -7454 408934
rect -7218 408698 480 408934
rect -8576 408676 480 408698
rect 583520 409254 592500 409276
rect 583520 409018 591142 409254
rect 591378 409018 592500 409254
rect 583520 408934 592500 409018
rect 583520 408698 591142 408934
rect 591378 408698 592500 408934
rect 583520 408676 592500 408698
rect -7636 408674 -7036 408676
rect 590960 408674 591560 408676
rect -5756 405676 -5156 405678
rect 589080 405676 589680 405678
rect -6696 405654 480 405676
rect -6696 405418 -5574 405654
rect -5338 405418 480 405654
rect -6696 405334 480 405418
rect -6696 405098 -5574 405334
rect -5338 405098 480 405334
rect -6696 405076 480 405098
rect 583520 405654 590620 405676
rect 583520 405418 589262 405654
rect 589498 405418 590620 405654
rect 583520 405334 590620 405418
rect 583520 405098 589262 405334
rect 589498 405098 590620 405334
rect 583520 405076 590620 405098
rect -5756 405074 -5156 405076
rect 589080 405074 589680 405076
rect -3876 402076 -3276 402078
rect 587200 402076 587800 402078
rect -4816 402054 480 402076
rect -4816 401818 -3694 402054
rect -3458 401818 480 402054
rect -4816 401734 480 401818
rect -4816 401498 -3694 401734
rect -3458 401498 480 401734
rect -4816 401476 480 401498
rect 583520 402054 588740 402076
rect 583520 401818 587382 402054
rect 587618 401818 588740 402054
rect 583520 401734 588740 401818
rect 583520 401498 587382 401734
rect 587618 401498 588740 401734
rect 583520 401476 588740 401498
rect -3876 401474 -3276 401476
rect 587200 401474 587800 401476
rect 545608 398480 546512 398486
rect -1996 398476 -1396 398478
rect 545608 398476 546546 398480
rect 585320 398476 585920 398478
rect -2936 398454 480 398476
rect -2936 398218 -1814 398454
rect -1578 398218 480 398454
rect -2936 398134 480 398218
rect -2936 397898 -1814 398134
rect -1578 397898 480 398134
rect -2936 397876 480 397898
rect 545608 398460 586860 398476
rect 545608 398224 545956 398460
rect 546192 398454 586860 398460
rect 546192 398224 585502 398454
rect 545608 398218 585502 398224
rect 585738 398218 586860 398454
rect 545608 398140 586860 398218
rect 545608 397904 545956 398140
rect 546192 398134 586860 398140
rect 546192 397904 585502 398134
rect 545608 397898 585502 397904
rect 585738 397898 586860 398134
rect 545608 397876 586860 397898
rect -1996 397874 -1396 397876
rect 585320 397874 585920 397876
rect -8576 391276 -7976 391278
rect 591900 391276 592500 391278
rect -8576 391254 480 391276
rect -8576 391018 -8394 391254
rect -8158 391018 480 391254
rect -8576 390934 480 391018
rect -8576 390698 -8394 390934
rect -8158 390698 480 390934
rect -8576 390676 480 390698
rect 583520 391254 592500 391276
rect 583520 391018 592082 391254
rect 592318 391018 592500 391254
rect 583520 390934 592500 391018
rect 583520 390698 592082 390934
rect 592318 390698 592500 390934
rect 583520 390676 592500 390698
rect -8576 390674 -7976 390676
rect 591900 390674 592500 390676
rect -6696 387676 -6096 387678
rect 590020 387676 590620 387678
rect -6696 387654 480 387676
rect -6696 387418 -6514 387654
rect -6278 387418 480 387654
rect -6696 387334 480 387418
rect -6696 387098 -6514 387334
rect -6278 387098 480 387334
rect -6696 387076 480 387098
rect 583520 387654 590620 387676
rect 583520 387418 590202 387654
rect 590438 387418 590620 387654
rect 583520 387334 590620 387418
rect 583520 387098 590202 387334
rect 590438 387098 590620 387334
rect 583520 387076 590620 387098
rect -6696 387074 -6096 387076
rect 590020 387074 590620 387076
rect -4816 384076 -4216 384078
rect 588140 384076 588740 384078
rect -4816 384054 480 384076
rect -4816 383818 -4634 384054
rect -4398 383818 480 384054
rect -4816 383734 480 383818
rect -4816 383498 -4634 383734
rect -4398 383498 480 383734
rect -4816 383476 480 383498
rect 583520 384054 588740 384076
rect 583520 383818 588322 384054
rect 588558 383818 588740 384054
rect 583520 383734 588740 383818
rect 583520 383498 588322 383734
rect 588558 383498 588740 383734
rect 583520 383476 588740 383498
rect -4816 383474 -4216 383476
rect 588140 383474 588740 383476
rect -2936 380476 -2336 380478
rect 586260 380476 586860 380478
rect -2936 380454 480 380476
rect -2936 380218 -2754 380454
rect -2518 380218 480 380454
rect -2936 380134 480 380218
rect -2936 379898 -2754 380134
rect -2518 379898 480 380134
rect -2936 379876 480 379898
rect 583500 380454 586860 380476
rect 583500 380218 586442 380454
rect 586678 380218 586860 380454
rect 583500 380134 586860 380218
rect 583500 379898 586442 380134
rect 586678 379898 586860 380134
rect 583500 379876 586860 379898
rect -2936 379874 -2336 379876
rect 586260 379874 586860 379876
rect -7636 373276 -7036 373278
rect 590960 373276 591560 373278
rect -8576 373254 480 373276
rect -8576 373018 -7454 373254
rect -7218 373018 480 373254
rect -8576 372934 480 373018
rect -8576 372698 -7454 372934
rect -7218 372698 480 372934
rect -8576 372676 480 372698
rect 583520 373254 592500 373276
rect 583520 373018 591142 373254
rect 591378 373018 592500 373254
rect 583520 372934 592500 373018
rect 583520 372698 591142 372934
rect 591378 372698 592500 372934
rect 583520 372676 592500 372698
rect -7636 372674 -7036 372676
rect 590960 372674 591560 372676
rect -5756 369676 -5156 369678
rect 589080 369676 589680 369678
rect -6696 369654 480 369676
rect -6696 369418 -5574 369654
rect -5338 369418 480 369654
rect -6696 369334 480 369418
rect -6696 369098 -5574 369334
rect -5338 369098 480 369334
rect -6696 369076 480 369098
rect 583520 369654 590620 369676
rect 583520 369418 589262 369654
rect 589498 369418 590620 369654
rect 583520 369334 590620 369418
rect 583520 369098 589262 369334
rect 589498 369098 590620 369334
rect 583520 369076 590620 369098
rect -5756 369074 -5156 369076
rect 589080 369074 589680 369076
rect -3876 366076 -3276 366078
rect 587200 366076 587800 366078
rect -4816 366054 480 366076
rect -4816 365818 -3694 366054
rect -3458 365818 480 366054
rect -4816 365734 480 365818
rect -4816 365498 -3694 365734
rect -3458 365498 480 365734
rect -4816 365476 480 365498
rect 583520 366054 588740 366076
rect 583520 365818 587382 366054
rect 587618 365818 588740 366054
rect 583520 365734 588740 365818
rect 583520 365498 587382 365734
rect 587618 365498 588740 365734
rect 583520 365476 588740 365498
rect -3876 365474 -3276 365476
rect 587200 365474 587800 365476
rect -1996 362476 -1396 362478
rect 585320 362476 585920 362478
rect -2936 362454 480 362476
rect -2936 362218 -1814 362454
rect -1578 362218 480 362454
rect -2936 362134 480 362218
rect -2936 361898 -1814 362134
rect -1578 361898 480 362134
rect -2936 361876 480 361898
rect 583520 362454 586860 362476
rect 583520 362218 585502 362454
rect 585738 362218 586860 362454
rect 583520 362134 586860 362218
rect 583520 361898 585502 362134
rect 585738 361898 586860 362134
rect 583520 361876 586860 361898
rect -1996 361874 -1396 361876
rect 585320 361874 585920 361876
rect -8576 355276 -7976 355278
rect 591900 355276 592500 355278
rect -8576 355254 480 355276
rect -8576 355018 -8394 355254
rect -8158 355018 480 355254
rect -8576 354934 480 355018
rect -8576 354698 -8394 354934
rect -8158 354698 480 354934
rect -8576 354676 480 354698
rect 583520 355254 592500 355276
rect 583520 355018 592082 355254
rect 592318 355018 592500 355254
rect 583520 354934 592500 355018
rect 583520 354698 592082 354934
rect 592318 354698 592500 354934
rect 583520 354676 592500 354698
rect -8576 354674 -7976 354676
rect 591900 354674 592500 354676
rect -6696 351676 -6096 351678
rect 590020 351676 590620 351678
rect -6696 351654 480 351676
rect -6696 351418 -6514 351654
rect -6278 351418 480 351654
rect -6696 351334 480 351418
rect -6696 351098 -6514 351334
rect -6278 351098 480 351334
rect -6696 351076 480 351098
rect 583520 351654 590620 351676
rect 583520 351418 590202 351654
rect 590438 351418 590620 351654
rect 583520 351334 590620 351418
rect 583520 351098 590202 351334
rect 590438 351098 590620 351334
rect 583520 351076 590620 351098
rect -6696 351074 -6096 351076
rect 590020 351074 590620 351076
rect -4816 348076 -4216 348078
rect 588140 348076 588740 348078
rect -4816 348054 480 348076
rect -4816 347818 -4634 348054
rect -4398 347818 480 348054
rect -4816 347734 480 347818
rect -4816 347498 -4634 347734
rect -4398 347498 480 347734
rect -4816 347476 480 347498
rect 583520 348054 588740 348076
rect 583520 347818 588322 348054
rect 588558 347818 588740 348054
rect 583520 347734 588740 347818
rect 583520 347498 588322 347734
rect 588558 347498 588740 347734
rect 583520 347476 588740 347498
rect -4816 347474 -4216 347476
rect 588140 347474 588740 347476
rect -2936 344476 -2336 344478
rect 586260 344476 586860 344478
rect -2936 344454 480 344476
rect -2936 344218 -2754 344454
rect -2518 344218 480 344454
rect -2936 344134 480 344218
rect -2936 343898 -2754 344134
rect -2518 343898 480 344134
rect -2936 343876 480 343898
rect 583520 344454 586860 344476
rect 583520 344218 586442 344454
rect 586678 344218 586860 344454
rect 583520 344134 586860 344218
rect 583520 343898 586442 344134
rect 586678 343898 586860 344134
rect 583520 343876 586860 343898
rect -2936 343874 -2336 343876
rect 586260 343874 586860 343876
rect -7636 337276 -7036 337278
rect 590960 337276 591560 337278
rect -8576 337254 480 337276
rect -8576 337018 -7454 337254
rect -7218 337018 480 337254
rect -8576 336934 480 337018
rect -8576 336698 -7454 336934
rect -7218 336698 480 336934
rect -8576 336676 480 336698
rect 583520 337254 592500 337276
rect 583520 337018 591142 337254
rect 591378 337018 592500 337254
rect 583520 336934 592500 337018
rect 583520 336698 591142 336934
rect 591378 336698 592500 336934
rect 583520 336676 592500 336698
rect -7636 336674 -7036 336676
rect 590960 336674 591560 336676
rect -5756 333676 -5156 333678
rect 589080 333676 589680 333678
rect -6696 333654 480 333676
rect -6696 333418 -5574 333654
rect -5338 333418 480 333654
rect -6696 333334 480 333418
rect -6696 333098 -5574 333334
rect -5338 333098 480 333334
rect -6696 333076 480 333098
rect 583520 333654 590620 333676
rect 583520 333418 589262 333654
rect 589498 333418 590620 333654
rect 583520 333334 590620 333418
rect 583520 333098 589262 333334
rect 589498 333098 590620 333334
rect 583520 333076 590620 333098
rect -5756 333074 -5156 333076
rect 589080 333074 589680 333076
rect -3876 330076 -3276 330078
rect 587200 330076 587800 330078
rect -4816 330054 480 330076
rect -4816 329818 -3694 330054
rect -3458 329818 480 330054
rect -4816 329734 480 329818
rect -4816 329498 -3694 329734
rect -3458 329498 480 329734
rect -4816 329476 480 329498
rect 583520 330054 588740 330076
rect 583520 329818 587382 330054
rect 587618 329818 588740 330054
rect 583520 329734 588740 329818
rect 583520 329498 587382 329734
rect 587618 329498 588740 329734
rect 583520 329476 588740 329498
rect -3876 329474 -3276 329476
rect 587200 329474 587800 329476
rect -1996 326476 -1396 326478
rect 585320 326476 585920 326478
rect -2936 326454 480 326476
rect -2936 326218 -1814 326454
rect -1578 326218 480 326454
rect -2936 326134 480 326218
rect -2936 325898 -1814 326134
rect -1578 325898 480 326134
rect -2936 325876 480 325898
rect 583520 326454 586860 326476
rect 583520 326218 585502 326454
rect 585738 326218 586860 326454
rect 583520 326134 586860 326218
rect 583520 325898 585502 326134
rect 585738 325898 586860 326134
rect 583520 325876 586860 325898
rect -1996 325874 -1396 325876
rect 585320 325874 585920 325876
rect -8576 319276 -7976 319278
rect 591900 319276 592500 319278
rect -8576 319254 480 319276
rect -8576 319018 -8394 319254
rect -8158 319018 480 319254
rect -8576 318934 480 319018
rect -8576 318698 -8394 318934
rect -8158 318698 480 318934
rect -8576 318676 480 318698
rect 583520 319254 592500 319276
rect 583520 319018 592082 319254
rect 592318 319018 592500 319254
rect 583520 318934 592500 319018
rect 583520 318698 592082 318934
rect 592318 318698 592500 318934
rect 583520 318676 592500 318698
rect -8576 318674 -7976 318676
rect 591900 318674 592500 318676
rect -6696 315676 -6096 315678
rect 590020 315676 590620 315678
rect -6696 315654 480 315676
rect -6696 315418 -6514 315654
rect -6278 315418 480 315654
rect -6696 315334 480 315418
rect -6696 315098 -6514 315334
rect -6278 315098 480 315334
rect -6696 315076 480 315098
rect 583520 315654 590620 315676
rect 583520 315418 590202 315654
rect 590438 315418 590620 315654
rect 583520 315334 590620 315418
rect 583520 315098 590202 315334
rect 590438 315098 590620 315334
rect 583520 315076 590620 315098
rect -6696 315074 -6096 315076
rect 590020 315074 590620 315076
rect -4816 312076 -4216 312078
rect 588140 312076 588740 312078
rect -4816 312054 480 312076
rect -4816 311818 -4634 312054
rect -4398 311818 480 312054
rect -4816 311734 480 311818
rect -4816 311498 -4634 311734
rect -4398 311498 480 311734
rect -4816 311476 480 311498
rect 583520 312054 588740 312076
rect 583520 311818 588322 312054
rect 588558 311818 588740 312054
rect 583520 311734 588740 311818
rect 583520 311498 588322 311734
rect 588558 311498 588740 311734
rect 583520 311476 588740 311498
rect -4816 311474 -4216 311476
rect 588140 311474 588740 311476
rect -2936 308476 -2336 308478
rect 586260 308476 586860 308478
rect -2936 308454 480 308476
rect -2936 308218 -2754 308454
rect -2518 308218 480 308454
rect -2936 308134 480 308218
rect -2936 307898 -2754 308134
rect -2518 307898 480 308134
rect -2936 307876 480 307898
rect 583520 308454 586860 308476
rect 583520 308218 586442 308454
rect 586678 308218 586860 308454
rect 583520 308134 586860 308218
rect 583520 307898 586442 308134
rect 586678 307898 586860 308134
rect 583520 307876 586860 307898
rect -2936 307874 -2336 307876
rect 586260 307874 586860 307876
rect -7636 301276 -7036 301278
rect 590960 301276 591560 301278
rect -8576 301254 480 301276
rect -8576 301018 -7454 301254
rect -7218 301018 480 301254
rect -8576 300934 480 301018
rect -8576 300698 -7454 300934
rect -7218 300698 480 300934
rect -8576 300676 480 300698
rect 583520 301254 592500 301276
rect 583520 301018 591142 301254
rect 591378 301018 592500 301254
rect 583520 300934 592500 301018
rect 583520 300698 591142 300934
rect 591378 300698 592500 300934
rect 583520 300676 592500 300698
rect -7636 300674 -7036 300676
rect 590960 300674 591560 300676
rect -5756 297676 -5156 297678
rect 589080 297676 589680 297678
rect -6696 297654 480 297676
rect -6696 297418 -5574 297654
rect -5338 297418 480 297654
rect -6696 297334 480 297418
rect -6696 297098 -5574 297334
rect -5338 297098 480 297334
rect -6696 297076 480 297098
rect 583520 297654 590620 297676
rect 583520 297418 589262 297654
rect 589498 297418 590620 297654
rect 583520 297334 590620 297418
rect 583520 297098 589262 297334
rect 589498 297098 590620 297334
rect 583520 297076 590620 297098
rect -5756 297074 -5156 297076
rect 589080 297074 589680 297076
rect -3876 294076 -3276 294078
rect 587200 294076 587800 294078
rect -4816 294054 480 294076
rect -4816 293818 -3694 294054
rect -3458 293818 480 294054
rect -4816 293734 480 293818
rect -4816 293498 -3694 293734
rect -3458 293498 480 293734
rect -4816 293476 480 293498
rect 583520 294054 588740 294076
rect 583520 293818 587382 294054
rect 587618 293818 588740 294054
rect 583520 293734 588740 293818
rect 583520 293498 587382 293734
rect 587618 293498 588740 293734
rect 583520 293476 588740 293498
rect -3876 293474 -3276 293476
rect 587200 293474 587800 293476
rect -1996 290476 -1396 290478
rect 585320 290476 585920 290478
rect -2936 290454 480 290476
rect -2936 290218 -1814 290454
rect -1578 290218 480 290454
rect -2936 290134 480 290218
rect -2936 289898 -1814 290134
rect -1578 289898 480 290134
rect -2936 289876 480 289898
rect 583520 290454 586860 290476
rect 583520 290218 585502 290454
rect 585738 290218 586860 290454
rect 583520 290134 586860 290218
rect 583520 289898 585502 290134
rect 585738 289898 586860 290134
rect 583520 289876 586860 289898
rect -1996 289874 -1396 289876
rect 585320 289874 585920 289876
rect -8576 283276 -7976 283278
rect 591900 283276 592500 283278
rect -8576 283254 480 283276
rect -8576 283018 -8394 283254
rect -8158 283018 480 283254
rect -8576 282934 480 283018
rect -8576 282698 -8394 282934
rect -8158 282698 480 282934
rect -8576 282676 480 282698
rect 583520 283254 592500 283276
rect 583520 283018 592082 283254
rect 592318 283018 592500 283254
rect 583520 282934 592500 283018
rect 583520 282698 592082 282934
rect 592318 282698 592500 282934
rect 583520 282676 592500 282698
rect -8576 282674 -7976 282676
rect 591900 282674 592500 282676
rect -6696 279676 -6096 279678
rect 590020 279676 590620 279678
rect -6696 279654 480 279676
rect -6696 279418 -6514 279654
rect -6278 279418 480 279654
rect -6696 279334 480 279418
rect -6696 279098 -6514 279334
rect -6278 279098 480 279334
rect -6696 279076 480 279098
rect 583520 279654 590620 279676
rect 583520 279418 590202 279654
rect 590438 279418 590620 279654
rect 583520 279334 590620 279418
rect 583520 279098 590202 279334
rect 590438 279098 590620 279334
rect 583520 279076 590620 279098
rect -6696 279074 -6096 279076
rect 590020 279074 590620 279076
rect -4816 276076 -4216 276078
rect 588140 276076 588740 276078
rect -4816 276054 480 276076
rect -4816 275818 -4634 276054
rect -4398 275818 480 276054
rect -4816 275734 480 275818
rect -4816 275498 -4634 275734
rect -4398 275498 480 275734
rect -4816 275476 480 275498
rect 583520 276054 588740 276076
rect 583520 275818 588322 276054
rect 588558 275818 588740 276054
rect 583520 275734 588740 275818
rect 583520 275498 588322 275734
rect 588558 275498 588740 275734
rect 583520 275476 588740 275498
rect -4816 275474 -4216 275476
rect 588140 275474 588740 275476
rect -2936 272476 -2336 272478
rect 586260 272476 586860 272478
rect -2936 272454 480 272476
rect -2936 272218 -2754 272454
rect -2518 272218 480 272454
rect -2936 272134 480 272218
rect -2936 271898 -2754 272134
rect -2518 271898 480 272134
rect -2936 271876 480 271898
rect 583520 272454 586860 272476
rect 583520 272218 586442 272454
rect 586678 272218 586860 272454
rect 583520 272134 586860 272218
rect 583520 271898 586442 272134
rect 586678 271898 586860 272134
rect 583520 271876 586860 271898
rect -2936 271874 -2336 271876
rect 586260 271874 586860 271876
rect -7636 265276 -7036 265278
rect 590960 265276 591560 265278
rect -8576 265254 480 265276
rect -8576 265018 -7454 265254
rect -7218 265018 480 265254
rect -8576 264934 480 265018
rect -8576 264698 -7454 264934
rect -7218 264698 480 264934
rect -8576 264676 480 264698
rect 583520 265254 592500 265276
rect 583520 265018 591142 265254
rect 591378 265018 592500 265254
rect 583520 264934 592500 265018
rect 583520 264698 591142 264934
rect 591378 264698 592500 264934
rect 583520 264676 592500 264698
rect -7636 264674 -7036 264676
rect 590960 264674 591560 264676
rect -5756 261676 -5156 261678
rect 589080 261676 589680 261678
rect -6696 261654 480 261676
rect -6696 261418 -5574 261654
rect -5338 261418 480 261654
rect -6696 261334 480 261418
rect -6696 261098 -5574 261334
rect -5338 261098 480 261334
rect -6696 261076 480 261098
rect 583520 261654 590620 261676
rect 583520 261418 589262 261654
rect 589498 261418 590620 261654
rect 583520 261334 590620 261418
rect 583520 261098 589262 261334
rect 589498 261098 590620 261334
rect 583520 261076 590620 261098
rect -5756 261074 -5156 261076
rect 589080 261074 589680 261076
rect -3876 258076 -3276 258078
rect 587200 258076 587800 258078
rect -4816 258054 480 258076
rect -4816 257818 -3694 258054
rect -3458 257818 480 258054
rect -4816 257734 480 257818
rect -4816 257498 -3694 257734
rect -3458 257498 480 257734
rect -4816 257476 480 257498
rect 583520 258054 588740 258076
rect 583520 257818 587382 258054
rect 587618 257818 588740 258054
rect 583520 257734 588740 257818
rect 583520 257498 587382 257734
rect 587618 257498 588740 257734
rect 583520 257476 588740 257498
rect -3876 257474 -3276 257476
rect 587200 257474 587800 257476
rect -1996 254476 -1396 254478
rect 585320 254476 585920 254478
rect -2936 254454 480 254476
rect -2936 254218 -1814 254454
rect -1578 254218 480 254454
rect -2936 254134 480 254218
rect -2936 253898 -1814 254134
rect -1578 253898 480 254134
rect -2936 253876 480 253898
rect 583520 254454 586860 254476
rect 583520 254218 585502 254454
rect 585738 254218 586860 254454
rect 583520 254134 586860 254218
rect 583520 253898 585502 254134
rect 585738 253898 586860 254134
rect 583520 253876 586860 253898
rect -1996 253874 -1396 253876
rect 585320 253874 585920 253876
rect -8576 247276 -7976 247278
rect 591900 247276 592500 247278
rect -8576 247254 480 247276
rect -8576 247018 -8394 247254
rect -8158 247018 480 247254
rect -8576 246934 480 247018
rect -8576 246698 -8394 246934
rect -8158 246698 480 246934
rect -8576 246676 480 246698
rect 583520 247254 592500 247276
rect 583520 247018 592082 247254
rect 592318 247018 592500 247254
rect 583520 246934 592500 247018
rect 583520 246698 592082 246934
rect 592318 246698 592500 246934
rect 583520 246676 592500 246698
rect -8576 246674 -7976 246676
rect 591900 246674 592500 246676
rect -6696 243676 -6096 243678
rect 590020 243676 590620 243678
rect -6696 243654 480 243676
rect -6696 243418 -6514 243654
rect -6278 243418 480 243654
rect -6696 243334 480 243418
rect -6696 243098 -6514 243334
rect -6278 243098 480 243334
rect -6696 243076 480 243098
rect 583520 243654 590620 243676
rect 583520 243418 590202 243654
rect 590438 243418 590620 243654
rect 583520 243334 590620 243418
rect 583520 243098 590202 243334
rect 590438 243098 590620 243334
rect 583520 243076 590620 243098
rect -6696 243074 -6096 243076
rect 590020 243074 590620 243076
rect -4816 240076 -4216 240078
rect 588140 240076 588740 240078
rect -4816 240054 480 240076
rect -4816 239818 -4634 240054
rect -4398 239818 480 240054
rect -4816 239734 480 239818
rect -4816 239498 -4634 239734
rect -4398 239498 480 239734
rect -4816 239476 480 239498
rect 583520 240054 588740 240076
rect 583520 239818 588322 240054
rect 588558 239818 588740 240054
rect 583520 239734 588740 239818
rect 583520 239498 588322 239734
rect 588558 239498 588740 239734
rect 583520 239476 588740 239498
rect -4816 239474 -4216 239476
rect 588140 239474 588740 239476
rect 544064 236480 544904 236484
rect -2936 236476 -2336 236478
rect 544016 236476 544930 236480
rect 586260 236476 586860 236478
rect -2936 236454 480 236476
rect -2936 236218 -2754 236454
rect -2518 236218 480 236454
rect -2936 236134 480 236218
rect -2936 235898 -2754 236134
rect -2518 235898 480 236134
rect -2936 235876 480 235898
rect 544016 236458 586860 236476
rect 544016 236222 544412 236458
rect 544648 236454 586860 236458
rect 544648 236222 586442 236454
rect 544016 236218 586442 236222
rect 586678 236218 586860 236454
rect 544016 236138 586860 236218
rect 544016 235902 544412 236138
rect 544648 236134 586860 236138
rect 544648 235902 586442 236134
rect 544016 235898 586442 235902
rect 586678 235898 586860 236134
rect 544016 235880 586860 235898
rect 544018 235876 586860 235880
rect -2936 235874 -2336 235876
rect 544064 235874 544904 235876
rect 586260 235874 586860 235876
rect -7636 229276 -7036 229278
rect 590960 229276 591560 229278
rect -8576 229254 480 229276
rect -8576 229018 -7454 229254
rect -7218 229018 480 229254
rect -8576 228934 480 229018
rect -8576 228698 -7454 228934
rect -7218 228698 480 228934
rect -8576 228676 480 228698
rect 583520 229254 592500 229276
rect 583520 229018 591142 229254
rect 591378 229018 592500 229254
rect 583520 228934 592500 229018
rect 583520 228698 591142 228934
rect 591378 228698 592500 228934
rect 583520 228676 592500 228698
rect -7636 228674 -7036 228676
rect 590960 228674 591560 228676
rect -5756 225676 -5156 225678
rect 589080 225676 589680 225678
rect -6696 225654 480 225676
rect -6696 225418 -5574 225654
rect -5338 225418 480 225654
rect -6696 225334 480 225418
rect -6696 225098 -5574 225334
rect -5338 225098 480 225334
rect -6696 225076 480 225098
rect 583520 225654 590620 225676
rect 583520 225418 589262 225654
rect 589498 225418 590620 225654
rect 583520 225334 590620 225418
rect 583520 225098 589262 225334
rect 589498 225098 590620 225334
rect 583520 225076 590620 225098
rect -5756 225074 -5156 225076
rect 589080 225074 589680 225076
rect -3876 222076 -3276 222078
rect 587200 222076 587800 222078
rect -4816 222054 480 222076
rect -4816 221818 -3694 222054
rect -3458 221818 480 222054
rect -4816 221734 480 221818
rect -4816 221498 -3694 221734
rect -3458 221498 480 221734
rect -4816 221476 480 221498
rect 583520 222054 588740 222076
rect 583520 221818 587382 222054
rect 587618 221818 588740 222054
rect 583520 221734 588740 221818
rect 583520 221498 587382 221734
rect 587618 221498 588740 221734
rect 583520 221476 588740 221498
rect -3876 221474 -3276 221476
rect 587200 221474 587800 221476
rect -1996 218476 -1396 218478
rect 585320 218476 585920 218478
rect -2936 218454 480 218476
rect -2936 218218 -1814 218454
rect -1578 218218 480 218454
rect -2936 218134 480 218218
rect -2936 217898 -1814 218134
rect -1578 217898 480 218134
rect -2936 217876 480 217898
rect 583520 218454 586860 218476
rect 583520 218218 585502 218454
rect 585738 218218 586860 218454
rect 583520 218134 586860 218218
rect 583520 217898 585502 218134
rect 585738 217898 586860 218134
rect 583520 217876 586860 217898
rect -1996 217874 -1396 217876
rect 585320 217874 585920 217876
rect -8576 211276 -7976 211278
rect 591900 211276 592500 211278
rect -8576 211254 480 211276
rect -8576 211018 -8394 211254
rect -8158 211018 480 211254
rect -8576 210934 480 211018
rect -8576 210698 -8394 210934
rect -8158 210698 480 210934
rect -8576 210676 480 210698
rect 583520 211254 592500 211276
rect 583520 211018 592082 211254
rect 592318 211018 592500 211254
rect 583520 210934 592500 211018
rect 583520 210698 592082 210934
rect 592318 210698 592500 210934
rect 583520 210676 592500 210698
rect -8576 210674 -7976 210676
rect 591900 210674 592500 210676
rect -6696 207676 -6096 207678
rect 590020 207676 590620 207678
rect -6696 207654 480 207676
rect -6696 207418 -6514 207654
rect -6278 207418 480 207654
rect -6696 207334 480 207418
rect -6696 207098 -6514 207334
rect -6278 207098 480 207334
rect -6696 207076 480 207098
rect 583520 207654 590620 207676
rect 583520 207418 590202 207654
rect 590438 207418 590620 207654
rect 583520 207334 590620 207418
rect 583520 207098 590202 207334
rect 590438 207098 590620 207334
rect 583520 207076 590620 207098
rect -6696 207074 -6096 207076
rect 590020 207074 590620 207076
rect -4816 204076 -4216 204078
rect 588140 204076 588740 204078
rect -4816 204054 480 204076
rect -4816 203818 -4634 204054
rect -4398 203818 480 204054
rect -4816 203734 480 203818
rect -4816 203498 -4634 203734
rect -4398 203498 480 203734
rect -4816 203476 480 203498
rect 583520 204054 588740 204076
rect 583520 203818 588322 204054
rect 588558 203818 588740 204054
rect 583520 203734 588740 203818
rect 583520 203498 588322 203734
rect 588558 203498 588740 203734
rect 583520 203476 588740 203498
rect -4816 203474 -4216 203476
rect 588140 203474 588740 203476
rect -2936 200476 -2336 200478
rect 586260 200476 586860 200478
rect -2936 200454 480 200476
rect -2936 200218 -2754 200454
rect -2518 200218 480 200454
rect -2936 200134 480 200218
rect -2936 199898 -2754 200134
rect -2518 199898 480 200134
rect -2936 199876 480 199898
rect 583520 200454 586860 200476
rect 583520 200218 586442 200454
rect 586678 200218 586860 200454
rect 583520 200134 586860 200218
rect 583520 199898 586442 200134
rect 586678 199898 586860 200134
rect 583520 199876 586860 199898
rect -2936 199874 -2336 199876
rect 586260 199874 586860 199876
rect -7636 193276 -7036 193278
rect 590960 193276 591560 193278
rect -8576 193254 480 193276
rect -8576 193018 -7454 193254
rect -7218 193018 480 193254
rect -8576 192934 480 193018
rect -8576 192698 -7454 192934
rect -7218 192698 480 192934
rect -8576 192676 480 192698
rect 583520 193254 592500 193276
rect 583520 193018 591142 193254
rect 591378 193018 592500 193254
rect 583520 192934 592500 193018
rect 583520 192698 591142 192934
rect 591378 192698 592500 192934
rect 583520 192676 592500 192698
rect -7636 192674 -7036 192676
rect 590960 192674 591560 192676
rect -5756 189676 -5156 189678
rect 589080 189676 589680 189678
rect -6696 189654 480 189676
rect -6696 189418 -5574 189654
rect -5338 189418 480 189654
rect -6696 189334 480 189418
rect -6696 189098 -5574 189334
rect -5338 189098 480 189334
rect -6696 189076 480 189098
rect 583520 189654 590620 189676
rect 583520 189418 589262 189654
rect 589498 189418 590620 189654
rect 583520 189334 590620 189418
rect 583520 189098 589262 189334
rect 589498 189098 590620 189334
rect 583520 189076 590620 189098
rect -5756 189074 -5156 189076
rect 589080 189074 589680 189076
rect -3876 186076 -3276 186078
rect 587200 186076 587800 186078
rect -4816 186054 480 186076
rect -4816 185818 -3694 186054
rect -3458 185818 480 186054
rect -4816 185734 480 185818
rect -4816 185498 -3694 185734
rect -3458 185498 480 185734
rect -4816 185476 480 185498
rect 583520 186054 588740 186076
rect 583520 185818 587382 186054
rect 587618 185818 588740 186054
rect 583520 185734 588740 185818
rect 583520 185498 587382 185734
rect 587618 185498 588740 185734
rect 583520 185476 588740 185498
rect -3876 185474 -3276 185476
rect 587200 185474 587800 185476
rect 544534 182490 545344 182494
rect 544534 182480 545444 182490
rect -1996 182476 -1396 182478
rect 544534 182476 545934 182480
rect 585320 182476 585920 182478
rect -2936 182454 480 182476
rect -2936 182218 -1814 182454
rect -1578 182218 480 182454
rect -2936 182134 480 182218
rect -2936 181898 -1814 182134
rect -1578 181898 480 182134
rect -2936 181876 480 181898
rect 544534 182468 586860 182476
rect 544534 182232 544876 182468
rect 545112 182454 586860 182468
rect 545112 182232 585502 182454
rect 544534 182218 585502 182232
rect 585738 182218 586860 182454
rect 544534 182148 586860 182218
rect 544534 181912 544876 182148
rect 545112 182134 586860 182148
rect 545112 181912 585502 182134
rect 544534 181898 585502 181912
rect 585738 181898 586860 182134
rect 544534 181876 586860 181898
rect -1996 181874 -1396 181876
rect 585320 181874 585920 181876
rect -8576 175276 -7976 175278
rect 591900 175276 592500 175278
rect -8576 175254 480 175276
rect -8576 175018 -8394 175254
rect -8158 175018 480 175254
rect -8576 174934 480 175018
rect -8576 174698 -8394 174934
rect -8158 174698 480 174934
rect -8576 174676 480 174698
rect 583520 175254 592500 175276
rect 583520 175018 592082 175254
rect 592318 175018 592500 175254
rect 583520 174934 592500 175018
rect 583520 174698 592082 174934
rect 592318 174698 592500 174934
rect 583520 174676 592500 174698
rect -8576 174674 -7976 174676
rect 591900 174674 592500 174676
rect -6696 171676 -6096 171678
rect 590020 171676 590620 171678
rect -6696 171654 480 171676
rect -6696 171418 -6514 171654
rect -6278 171418 480 171654
rect -6696 171334 480 171418
rect -6696 171098 -6514 171334
rect -6278 171098 480 171334
rect -6696 171076 480 171098
rect 583520 171654 590620 171676
rect 583520 171418 590202 171654
rect 590438 171418 590620 171654
rect 583520 171334 590620 171418
rect 583520 171098 590202 171334
rect 590438 171098 590620 171334
rect 583520 171076 590620 171098
rect -6696 171074 -6096 171076
rect 590020 171074 590620 171076
rect -4816 168076 -4216 168078
rect 588140 168076 588740 168078
rect -4816 168054 480 168076
rect -4816 167818 -4634 168054
rect -4398 167818 480 168054
rect -4816 167734 480 167818
rect -4816 167498 -4634 167734
rect -4398 167498 480 167734
rect -4816 167476 480 167498
rect 583520 168054 588740 168076
rect 583520 167818 588322 168054
rect 588558 167818 588740 168054
rect 583520 167734 588740 167818
rect 583520 167498 588322 167734
rect 588558 167498 588740 167734
rect 583520 167476 588740 167498
rect -4816 167474 -4216 167476
rect 588140 167474 588740 167476
rect -2936 164476 -2336 164478
rect 586260 164476 586860 164478
rect -2936 164454 480 164476
rect -2936 164218 -2754 164454
rect -2518 164218 480 164454
rect -2936 164134 480 164218
rect -2936 163898 -2754 164134
rect -2518 163898 480 164134
rect -2936 163876 480 163898
rect 583520 164454 586860 164476
rect 583520 164218 586442 164454
rect 586678 164218 586860 164454
rect 583520 164134 586860 164218
rect 583520 163898 586442 164134
rect 586678 163898 586860 164134
rect 583520 163876 586860 163898
rect -2936 163874 -2336 163876
rect 586260 163874 586860 163876
rect -7636 157276 -7036 157278
rect 590960 157276 591560 157278
rect -8576 157254 480 157276
rect -8576 157018 -7454 157254
rect -7218 157018 480 157254
rect -8576 156934 480 157018
rect -8576 156698 -7454 156934
rect -7218 156698 480 156934
rect -8576 156676 480 156698
rect 583520 157254 592500 157276
rect 583520 157018 591142 157254
rect 591378 157018 592500 157254
rect 583520 156934 592500 157018
rect 583520 156698 591142 156934
rect 591378 156698 592500 156934
rect 583520 156676 592500 156698
rect -7636 156674 -7036 156676
rect 590960 156674 591560 156676
rect -5756 153676 -5156 153678
rect 589080 153676 589680 153678
rect -6696 153654 480 153676
rect -6696 153418 -5574 153654
rect -5338 153418 480 153654
rect -6696 153334 480 153418
rect -6696 153098 -5574 153334
rect -5338 153098 480 153334
rect -6696 153076 480 153098
rect 583520 153654 590620 153676
rect 583520 153418 589262 153654
rect 589498 153418 590620 153654
rect 583520 153334 590620 153418
rect 583520 153098 589262 153334
rect 589498 153098 590620 153334
rect 583520 153076 590620 153098
rect -5756 153074 -5156 153076
rect 589080 153074 589680 153076
rect -3876 150076 -3276 150078
rect 587200 150076 587800 150078
rect -4816 150054 480 150076
rect -4816 149818 -3694 150054
rect -3458 149818 480 150054
rect -4816 149734 480 149818
rect -4816 149498 -3694 149734
rect -3458 149498 480 149734
rect -4816 149476 480 149498
rect 583520 150054 588740 150076
rect 583520 149818 587382 150054
rect 587618 149818 588740 150054
rect 583520 149734 588740 149818
rect 583520 149498 587382 149734
rect 587618 149498 588740 149734
rect 583520 149476 588740 149498
rect -3876 149474 -3276 149476
rect 587200 149474 587800 149476
rect -1996 146476 -1396 146478
rect 585320 146476 585920 146478
rect -2936 146454 480 146476
rect -2936 146218 -1814 146454
rect -1578 146218 480 146454
rect -2936 146134 480 146218
rect -2936 145898 -1814 146134
rect -1578 145898 480 146134
rect -2936 145876 480 145898
rect 583520 146454 586860 146476
rect 583520 146218 585502 146454
rect 585738 146218 586860 146454
rect 583520 146134 586860 146218
rect 583520 145898 585502 146134
rect 585738 145898 586860 146134
rect 583520 145876 586860 145898
rect -1996 145874 -1396 145876
rect 585320 145874 585920 145876
rect -8576 139276 -7976 139278
rect 591900 139276 592500 139278
rect -8576 139254 480 139276
rect -8576 139018 -8394 139254
rect -8158 139018 480 139254
rect -8576 138934 480 139018
rect -8576 138698 -8394 138934
rect -8158 138698 480 138934
rect -8576 138676 480 138698
rect 583520 139254 592500 139276
rect 583520 139018 592082 139254
rect 592318 139018 592500 139254
rect 583520 138934 592500 139018
rect 583520 138698 592082 138934
rect 592318 138698 592500 138934
rect 583520 138676 592500 138698
rect -8576 138674 -7976 138676
rect 591900 138674 592500 138676
rect -6696 135676 -6096 135678
rect 590020 135676 590620 135678
rect -6696 135654 480 135676
rect -6696 135418 -6514 135654
rect -6278 135418 480 135654
rect -6696 135334 480 135418
rect -6696 135098 -6514 135334
rect -6278 135098 480 135334
rect -6696 135076 480 135098
rect 583520 135654 590620 135676
rect 583520 135418 590202 135654
rect 590438 135418 590620 135654
rect 583520 135334 590620 135418
rect 583520 135098 590202 135334
rect 590438 135098 590620 135334
rect 583520 135076 590620 135098
rect -6696 135074 -6096 135076
rect 590020 135074 590620 135076
rect -4816 132076 -4216 132078
rect 588140 132076 588740 132078
rect -4816 132054 480 132076
rect -4816 131818 -4634 132054
rect -4398 131818 480 132054
rect -4816 131734 480 131818
rect -4816 131498 -4634 131734
rect -4398 131498 480 131734
rect -4816 131476 480 131498
rect 583520 132054 588740 132076
rect 583520 131818 588322 132054
rect 588558 131818 588740 132054
rect 583520 131734 588740 131818
rect 583520 131498 588322 131734
rect 588558 131498 588740 131734
rect 583520 131476 588740 131498
rect -4816 131474 -4216 131476
rect 588140 131474 588740 131476
rect -2936 128476 -2336 128478
rect 586260 128476 586860 128478
rect -2936 128454 480 128476
rect -2936 128218 -2754 128454
rect -2518 128218 480 128454
rect -2936 128134 480 128218
rect -2936 127898 -2754 128134
rect -2518 127898 480 128134
rect -2936 127876 480 127898
rect 583520 128454 586860 128476
rect 583520 128218 586442 128454
rect 586678 128218 586860 128454
rect 583520 128134 586860 128218
rect 583520 127898 586442 128134
rect 586678 127898 586860 128134
rect 583520 127876 586860 127898
rect -2936 127874 -2336 127876
rect 586260 127874 586860 127876
rect -7636 121276 -7036 121278
rect 590960 121276 591560 121278
rect -8576 121254 480 121276
rect -8576 121018 -7454 121254
rect -7218 121018 480 121254
rect -8576 120934 480 121018
rect -8576 120698 -7454 120934
rect -7218 120698 480 120934
rect -8576 120676 480 120698
rect 583520 121254 592500 121276
rect 583520 121018 591142 121254
rect 591378 121018 592500 121254
rect 583520 120934 592500 121018
rect 583520 120698 591142 120934
rect 591378 120698 592500 120934
rect 583520 120676 592500 120698
rect -7636 120674 -7036 120676
rect 590960 120674 591560 120676
rect -5756 117676 -5156 117678
rect 589080 117676 589680 117678
rect -6696 117654 480 117676
rect -6696 117418 -5574 117654
rect -5338 117418 480 117654
rect -6696 117334 480 117418
rect -6696 117098 -5574 117334
rect -5338 117098 480 117334
rect -6696 117076 480 117098
rect 583520 117654 590620 117676
rect 583520 117418 589262 117654
rect 589498 117418 590620 117654
rect 583520 117334 590620 117418
rect 583520 117098 589262 117334
rect 589498 117098 590620 117334
rect 583520 117076 590620 117098
rect -5756 117074 -5156 117076
rect 589080 117074 589680 117076
rect -3876 114076 -3276 114078
rect 587200 114076 587800 114078
rect -4816 114054 480 114076
rect -4816 113818 -3694 114054
rect -3458 113818 480 114054
rect -4816 113734 480 113818
rect -4816 113498 -3694 113734
rect -3458 113498 480 113734
rect -4816 113476 480 113498
rect 583520 114054 588740 114076
rect 583520 113818 587382 114054
rect 587618 113818 588740 114054
rect 583520 113734 588740 113818
rect 583520 113498 587382 113734
rect 587618 113498 588740 113734
rect 583520 113476 588740 113498
rect -3876 113474 -3276 113476
rect 587200 113474 587800 113476
rect -1996 110476 -1396 110478
rect 585320 110476 585920 110478
rect -2936 110454 480 110476
rect -2936 110218 -1814 110454
rect -1578 110218 480 110454
rect -2936 110134 480 110218
rect -2936 109898 -1814 110134
rect -1578 109898 480 110134
rect -2936 109876 480 109898
rect 583520 110454 586860 110476
rect 583520 110218 585502 110454
rect 585738 110218 586860 110454
rect 583520 110134 586860 110218
rect 583520 109898 585502 110134
rect 585738 109898 586860 110134
rect 583520 109876 586860 109898
rect -1996 109874 -1396 109876
rect 585320 109874 585920 109876
rect -8576 103276 -7976 103278
rect 591900 103276 592500 103278
rect -8576 103254 480 103276
rect -8576 103018 -8394 103254
rect -8158 103018 480 103254
rect -8576 102934 480 103018
rect -8576 102698 -8394 102934
rect -8158 102698 480 102934
rect -8576 102676 480 102698
rect 583520 103254 592500 103276
rect 583520 103018 592082 103254
rect 592318 103018 592500 103254
rect 583520 102934 592500 103018
rect 583520 102698 592082 102934
rect 592318 102698 592500 102934
rect 583520 102676 592500 102698
rect -8576 102674 -7976 102676
rect 591900 102674 592500 102676
rect -6696 99676 -6096 99678
rect 590020 99676 590620 99678
rect -6696 99654 480 99676
rect -6696 99418 -6514 99654
rect -6278 99418 480 99654
rect -6696 99334 480 99418
rect -6696 99098 -6514 99334
rect -6278 99098 480 99334
rect -6696 99076 480 99098
rect 583520 99654 590620 99676
rect 583520 99418 590202 99654
rect 590438 99418 590620 99654
rect 583520 99334 590620 99418
rect 583520 99098 590202 99334
rect 590438 99098 590620 99334
rect 583520 99076 590620 99098
rect -6696 99074 -6096 99076
rect 590020 99074 590620 99076
rect -4816 96076 -4216 96078
rect 588140 96076 588740 96078
rect -4816 96054 480 96076
rect -4816 95818 -4634 96054
rect -4398 95818 480 96054
rect -4816 95734 480 95818
rect -4816 95498 -4634 95734
rect -4398 95498 480 95734
rect -4816 95476 480 95498
rect 583520 96054 588740 96076
rect 583520 95818 588322 96054
rect 588558 95818 588740 96054
rect 583520 95734 588740 95818
rect 583520 95498 588322 95734
rect 588558 95498 588740 95734
rect 583520 95476 588740 95498
rect -4816 95474 -4216 95476
rect 588140 95474 588740 95476
rect -2936 92476 -2336 92478
rect 586260 92476 586860 92478
rect -2936 92454 480 92476
rect -2936 92218 -2754 92454
rect -2518 92218 480 92454
rect -2936 92134 480 92218
rect -2936 91898 -2754 92134
rect -2518 91898 480 92134
rect -2936 91876 480 91898
rect 583520 92454 586860 92476
rect 583520 92218 586442 92454
rect 586678 92218 586860 92454
rect 583520 92134 586860 92218
rect 583520 91898 586442 92134
rect 586678 91898 586860 92134
rect 583520 91876 586860 91898
rect -2936 91874 -2336 91876
rect 586260 91874 586860 91876
rect -7636 85276 -7036 85278
rect 590960 85276 591560 85278
rect -8576 85254 480 85276
rect -8576 85018 -7454 85254
rect -7218 85018 480 85254
rect -8576 84934 480 85018
rect -8576 84698 -7454 84934
rect -7218 84698 480 84934
rect -8576 84676 480 84698
rect 583520 85254 592500 85276
rect 583520 85018 591142 85254
rect 591378 85018 592500 85254
rect 583520 84934 592500 85018
rect 583520 84698 591142 84934
rect 591378 84698 592500 84934
rect 583520 84676 592500 84698
rect -7636 84674 -7036 84676
rect 590960 84674 591560 84676
rect -5756 81676 -5156 81678
rect 589080 81676 589680 81678
rect -6696 81654 480 81676
rect -6696 81418 -5574 81654
rect -5338 81418 480 81654
rect -6696 81334 480 81418
rect -6696 81098 -5574 81334
rect -5338 81098 480 81334
rect -6696 81076 480 81098
rect 583520 81654 590620 81676
rect 583520 81418 589262 81654
rect 589498 81418 590620 81654
rect 583520 81334 590620 81418
rect 583520 81098 589262 81334
rect 589498 81098 590620 81334
rect 583520 81076 590620 81098
rect -5756 81074 -5156 81076
rect 589080 81074 589680 81076
rect -3876 78076 -3276 78078
rect 587200 78076 587800 78078
rect -4816 78054 480 78076
rect -4816 77818 -3694 78054
rect -3458 77818 480 78054
rect -4816 77734 480 77818
rect -4816 77498 -3694 77734
rect -3458 77498 480 77734
rect -4816 77476 480 77498
rect 583520 78054 588740 78076
rect 583520 77818 587382 78054
rect 587618 77818 588740 78054
rect 583520 77734 588740 77818
rect 583520 77498 587382 77734
rect 587618 77498 588740 77734
rect 583520 77476 588740 77498
rect -3876 77474 -3276 77476
rect 587200 77474 587800 77476
rect -1996 74476 -1396 74478
rect 585320 74476 585920 74478
rect -2936 74454 480 74476
rect -2936 74218 -1814 74454
rect -1578 74218 480 74454
rect -2936 74134 480 74218
rect -2936 73898 -1814 74134
rect -1578 73898 480 74134
rect -2936 73876 480 73898
rect 583520 74454 586860 74476
rect 583520 74218 585502 74454
rect 585738 74218 586860 74454
rect 583520 74134 586860 74218
rect 583520 73898 585502 74134
rect 585738 73898 586860 74134
rect 583520 73876 586860 73898
rect -1996 73874 -1396 73876
rect 585320 73874 585920 73876
rect -8576 67276 -7976 67278
rect 591900 67276 592500 67278
rect -8576 67254 480 67276
rect -8576 67018 -8394 67254
rect -8158 67018 480 67254
rect -8576 66934 480 67018
rect -8576 66698 -8394 66934
rect -8158 66698 480 66934
rect -8576 66676 480 66698
rect 583520 67254 592500 67276
rect 583520 67018 592082 67254
rect 592318 67018 592500 67254
rect 583520 66934 592500 67018
rect 583520 66698 592082 66934
rect 592318 66698 592500 66934
rect 583520 66676 592500 66698
rect -8576 66674 -7976 66676
rect 591900 66674 592500 66676
rect -6696 63676 -6096 63678
rect 590020 63676 590620 63678
rect -6696 63654 480 63676
rect -6696 63418 -6514 63654
rect -6278 63418 480 63654
rect -6696 63334 480 63418
rect -6696 63098 -6514 63334
rect -6278 63098 480 63334
rect -6696 63076 480 63098
rect 583520 63654 590620 63676
rect 583520 63418 590202 63654
rect 590438 63418 590620 63654
rect 583520 63334 590620 63418
rect 583520 63098 590202 63334
rect 590438 63098 590620 63334
rect 583520 63076 590620 63098
rect -6696 63074 -6096 63076
rect 590020 63074 590620 63076
rect -4816 60076 -4216 60078
rect 588140 60076 588740 60078
rect -4816 60054 480 60076
rect -4816 59818 -4634 60054
rect -4398 59818 480 60054
rect -4816 59734 480 59818
rect -4816 59498 -4634 59734
rect -4398 59498 480 59734
rect -4816 59476 480 59498
rect 583520 60054 588740 60076
rect 583520 59818 588322 60054
rect 588558 59818 588740 60054
rect 583520 59734 588740 59818
rect 583520 59498 588322 59734
rect 588558 59498 588740 59734
rect 583520 59476 588740 59498
rect -4816 59474 -4216 59476
rect 588140 59474 588740 59476
rect -2936 56476 -2336 56478
rect 586260 56476 586860 56478
rect -2936 56454 480 56476
rect -2936 56218 -2754 56454
rect -2518 56218 480 56454
rect -2936 56134 480 56218
rect -2936 55898 -2754 56134
rect -2518 55898 480 56134
rect -2936 55876 480 55898
rect 583520 56454 586860 56476
rect 583520 56218 586442 56454
rect 586678 56218 586860 56454
rect 583520 56134 586860 56218
rect 583520 55898 586442 56134
rect 586678 55898 586860 56134
rect 583520 55876 586860 55898
rect -2936 55874 -2336 55876
rect 586260 55874 586860 55876
rect -7636 49276 -7036 49278
rect 590960 49276 591560 49278
rect -8576 49254 480 49276
rect -8576 49018 -7454 49254
rect -7218 49018 480 49254
rect -8576 48934 480 49018
rect -8576 48698 -7454 48934
rect -7218 48698 480 48934
rect -8576 48676 480 48698
rect 583520 49254 592500 49276
rect 583520 49018 591142 49254
rect 591378 49018 592500 49254
rect 583520 48934 592500 49018
rect 583520 48698 591142 48934
rect 591378 48698 592500 48934
rect 583520 48676 592500 48698
rect -7636 48674 -7036 48676
rect 590960 48674 591560 48676
rect -5756 45676 -5156 45678
rect 589080 45676 589680 45678
rect -6696 45654 480 45676
rect -6696 45418 -5574 45654
rect -5338 45418 480 45654
rect -6696 45334 480 45418
rect -6696 45098 -5574 45334
rect -5338 45098 480 45334
rect -6696 45076 480 45098
rect 583520 45654 590620 45676
rect 583520 45418 589262 45654
rect 589498 45418 590620 45654
rect 583520 45334 590620 45418
rect 583520 45098 589262 45334
rect 589498 45098 590620 45334
rect 583520 45076 590620 45098
rect -5756 45074 -5156 45076
rect 589080 45074 589680 45076
rect -3876 42076 -3276 42078
rect 587200 42076 587800 42078
rect -4816 42054 480 42076
rect -4816 41818 -3694 42054
rect -3458 41818 480 42054
rect -4816 41734 480 41818
rect -4816 41498 -3694 41734
rect -3458 41498 480 41734
rect -4816 41476 480 41498
rect 583520 42054 588740 42076
rect 583520 41818 587382 42054
rect 587618 41818 588740 42054
rect 583520 41734 588740 41818
rect 583520 41498 587382 41734
rect 587618 41498 588740 41734
rect 583520 41476 588740 41498
rect -3876 41474 -3276 41476
rect 587200 41474 587800 41476
rect -1996 38476 -1396 38478
rect 585320 38476 585920 38478
rect -2936 38454 480 38476
rect -2936 38218 -1814 38454
rect -1578 38218 480 38454
rect -2936 38134 480 38218
rect -2936 37898 -1814 38134
rect -1578 37898 480 38134
rect -2936 37876 480 37898
rect 583520 38454 586860 38476
rect 583520 38218 585502 38454
rect 585738 38218 586860 38454
rect 583520 38134 586860 38218
rect 583520 37898 585502 38134
rect 585738 37898 586860 38134
rect 583520 37876 586860 37898
rect -1996 37874 -1396 37876
rect 585320 37874 585920 37876
rect -8576 31276 -7976 31278
rect 591900 31276 592500 31278
rect -8576 31254 480 31276
rect -8576 31018 -8394 31254
rect -8158 31018 480 31254
rect -8576 30934 480 31018
rect -8576 30698 -8394 30934
rect -8158 30698 480 30934
rect -8576 30676 480 30698
rect 583520 31254 592500 31276
rect 583520 31018 592082 31254
rect 592318 31018 592500 31254
rect 583520 30934 592500 31018
rect 583520 30698 592082 30934
rect 592318 30698 592500 30934
rect 583520 30676 592500 30698
rect -8576 30674 -7976 30676
rect 591900 30674 592500 30676
rect -6696 27676 -6096 27678
rect 590020 27676 590620 27678
rect -6696 27654 480 27676
rect -6696 27418 -6514 27654
rect -6278 27418 480 27654
rect -6696 27334 480 27418
rect -6696 27098 -6514 27334
rect -6278 27098 480 27334
rect -6696 27076 480 27098
rect 583520 27654 590620 27676
rect 583520 27418 590202 27654
rect 590438 27418 590620 27654
rect 583520 27334 590620 27418
rect 583520 27098 590202 27334
rect 590438 27098 590620 27334
rect 583520 27076 590620 27098
rect -6696 27074 -6096 27076
rect 590020 27074 590620 27076
rect -4816 24076 -4216 24078
rect 588140 24076 588740 24078
rect -4816 24054 480 24076
rect -4816 23818 -4634 24054
rect -4398 23818 480 24054
rect -4816 23734 480 23818
rect -4816 23498 -4634 23734
rect -4398 23498 480 23734
rect -4816 23476 480 23498
rect 583520 24054 588740 24076
rect 583520 23818 588322 24054
rect 588558 23818 588740 24054
rect 583520 23734 588740 23818
rect 583520 23498 588322 23734
rect 588558 23498 588740 23734
rect 583520 23476 588740 23498
rect -4816 23474 -4216 23476
rect 588140 23474 588740 23476
rect -2936 20476 -2336 20478
rect 586260 20476 586860 20478
rect -2936 20454 480 20476
rect -2936 20218 -2754 20454
rect -2518 20218 480 20454
rect -2936 20134 480 20218
rect -2936 19898 -2754 20134
rect -2518 19898 480 20134
rect -2936 19876 480 19898
rect 583520 20454 586860 20476
rect 583520 20218 586442 20454
rect 586678 20218 586860 20454
rect 583520 20134 586860 20218
rect 583520 19898 586442 20134
rect 586678 19898 586860 20134
rect 583520 19876 586860 19898
rect -2936 19874 -2336 19876
rect 586260 19874 586860 19876
rect -7636 13276 -7036 13278
rect 590960 13276 591560 13278
rect -8576 13254 480 13276
rect -8576 13018 -7454 13254
rect -7218 13018 480 13254
rect -8576 12934 480 13018
rect -8576 12698 -7454 12934
rect -7218 12698 480 12934
rect -8576 12676 480 12698
rect 583520 13254 592500 13276
rect 583520 13018 591142 13254
rect 591378 13018 592500 13254
rect 583520 12934 592500 13018
rect 583520 12698 591142 12934
rect 591378 12698 592500 12934
rect 583520 12676 592500 12698
rect -7636 12674 -7036 12676
rect 590960 12674 591560 12676
rect -5756 9676 -5156 9678
rect 589080 9676 589680 9678
rect -6696 9654 480 9676
rect -6696 9418 -5574 9654
rect -5338 9418 480 9654
rect -6696 9334 480 9418
rect -6696 9098 -5574 9334
rect -5338 9098 480 9334
rect -6696 9076 480 9098
rect 583520 9654 590620 9676
rect 583520 9418 589262 9654
rect 589498 9418 590620 9654
rect 583520 9334 590620 9418
rect 583520 9098 589262 9334
rect 589498 9098 590620 9334
rect 583520 9076 590620 9098
rect -5756 9074 -5156 9076
rect 589080 9074 589680 9076
rect -3876 6076 -3276 6078
rect 587200 6076 587800 6078
rect -4816 6054 480 6076
rect -4816 5818 -3694 6054
rect -3458 5818 480 6054
rect -4816 5734 480 5818
rect -4816 5498 -3694 5734
rect -3458 5498 480 5734
rect -4816 5476 480 5498
rect 583520 6054 588740 6076
rect 583520 5818 587382 6054
rect 587618 5818 588740 6054
rect 583520 5734 588740 5818
rect 583520 5498 587382 5734
rect 587618 5498 588740 5734
rect 583520 5476 588740 5498
rect -3876 5474 -3276 5476
rect 587200 5474 587800 5476
rect -1996 2476 -1396 2478
rect 585320 2476 585920 2478
rect -2936 2454 480 2476
rect -2936 2218 -1814 2454
rect -1578 2218 480 2454
rect -2936 2134 480 2218
rect -2936 1898 -1814 2134
rect -1578 1898 480 2134
rect -2936 1876 480 1898
rect 583520 2454 586860 2476
rect 583520 2218 585502 2454
rect 585738 2218 586860 2454
rect 583520 2134 586860 2218
rect 583520 1898 585502 2134
rect 585738 1898 586860 2134
rect 583520 1876 586860 1898
rect -1996 1874 -1396 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 148404 -2204 149004 -2202
rect 184404 -2204 185004 -2202
rect 220404 -2204 221004 -2202
rect 256404 -2204 257004 -2202
rect 292404 -2204 293004 -2202
rect 328404 -2204 329004 -2202
rect 364404 -2204 365004 -2202
rect 400404 -2204 401004 -2202
rect 436404 -2204 437004 -2202
rect 472404 -2204 473004 -2202
rect 508404 -2204 509004 -2202
rect 544404 -2204 545004 -2202
rect 580404 -2204 581004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 4586 -2226
rect 4822 -2462 40586 -2226
rect 40822 -2462 76586 -2226
rect 76822 -2462 112586 -2226
rect 112822 -2462 148586 -2226
rect 148822 -2462 184586 -2226
rect 184822 -2462 220586 -2226
rect 220822 -2462 256586 -2226
rect 256822 -2462 292586 -2226
rect 292822 -2462 328586 -2226
rect 328822 -2462 364586 -2226
rect 364822 -2462 400586 -2226
rect 400822 -2462 436586 -2226
rect 436822 -2462 472586 -2226
rect 472822 -2462 508586 -2226
rect 508822 -2462 544586 -2226
rect 544822 -2462 580586 -2226
rect 580822 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 4586 -2546
rect 4822 -2782 40586 -2546
rect 40822 -2782 76586 -2546
rect 76822 -2782 112586 -2546
rect 112822 -2782 148586 -2546
rect 148822 -2782 184586 -2546
rect 184822 -2782 220586 -2546
rect 220822 -2782 256586 -2546
rect 256822 -2782 292586 -2546
rect 292822 -2782 328586 -2546
rect 328822 -2782 364586 -2546
rect 364822 -2782 400586 -2546
rect 400822 -2782 436586 -2546
rect 436822 -2782 472586 -2546
rect 472822 -2782 508586 -2546
rect 508822 -2782 544586 -2546
rect 544822 -2782 580586 -2546
rect 580822 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 148404 -2806 149004 -2804
rect 184404 -2806 185004 -2804
rect 220404 -2806 221004 -2804
rect 256404 -2806 257004 -2804
rect 292404 -2806 293004 -2804
rect 328404 -2806 329004 -2804
rect 364404 -2806 365004 -2804
rect 400404 -2806 401004 -2804
rect 436404 -2806 437004 -2804
rect 472404 -2806 473004 -2804
rect 508404 -2806 509004 -2804
rect 544404 -2806 545004 -2804
rect 580404 -2806 581004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 130404 -3144 131004 -3142
rect 166404 -3144 167004 -3142
rect 202404 -3144 203004 -3142
rect 238404 -3144 239004 -3142
rect 274404 -3144 275004 -3142
rect 310404 -3144 311004 -3142
rect 346404 -3144 347004 -3142
rect 382404 -3144 383004 -3142
rect 418404 -3144 419004 -3142
rect 454404 -3144 455004 -3142
rect 490404 -3144 491004 -3142
rect 526404 -3144 527004 -3142
rect 562404 -3144 563004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 22586 -3166
rect 22822 -3402 58586 -3166
rect 58822 -3402 94586 -3166
rect 94822 -3402 130586 -3166
rect 130822 -3402 166586 -3166
rect 166822 -3402 202586 -3166
rect 202822 -3402 238586 -3166
rect 238822 -3402 274586 -3166
rect 274822 -3402 310586 -3166
rect 310822 -3402 346586 -3166
rect 346822 -3402 382586 -3166
rect 382822 -3402 418586 -3166
rect 418822 -3402 454586 -3166
rect 454822 -3402 490586 -3166
rect 490822 -3402 526586 -3166
rect 526822 -3402 562586 -3166
rect 562822 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 22586 -3486
rect 22822 -3722 58586 -3486
rect 58822 -3722 94586 -3486
rect 94822 -3722 130586 -3486
rect 130822 -3722 166586 -3486
rect 166822 -3722 202586 -3486
rect 202822 -3722 238586 -3486
rect 238822 -3722 274586 -3486
rect 274822 -3722 310586 -3486
rect 310822 -3722 346586 -3486
rect 346822 -3722 382586 -3486
rect 382822 -3722 418586 -3486
rect 418822 -3722 454586 -3486
rect 454822 -3722 490586 -3486
rect 490822 -3722 526586 -3486
rect 526822 -3722 562586 -3486
rect 562822 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 130404 -3746 131004 -3744
rect 166404 -3746 167004 -3744
rect 202404 -3746 203004 -3744
rect 238404 -3746 239004 -3744
rect 274404 -3746 275004 -3744
rect 310404 -3746 311004 -3744
rect 346404 -3746 347004 -3744
rect 382404 -3746 383004 -3744
rect 418404 -3746 419004 -3744
rect 454404 -3746 455004 -3744
rect 490404 -3746 491004 -3744
rect 526404 -3746 527004 -3744
rect 562404 -3746 563004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 152004 -4084 152604 -4082
rect 188004 -4084 188604 -4082
rect 224004 -4084 224604 -4082
rect 260004 -4084 260604 -4082
rect 296004 -4084 296604 -4082
rect 332004 -4084 332604 -4082
rect 368004 -4084 368604 -4082
rect 404004 -4084 404604 -4082
rect 440004 -4084 440604 -4082
rect 476004 -4084 476604 -4082
rect 512004 -4084 512604 -4082
rect 548004 -4084 548604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 8186 -4106
rect 8422 -4342 44186 -4106
rect 44422 -4342 80186 -4106
rect 80422 -4342 116186 -4106
rect 116422 -4342 152186 -4106
rect 152422 -4342 188186 -4106
rect 188422 -4342 224186 -4106
rect 224422 -4342 260186 -4106
rect 260422 -4342 296186 -4106
rect 296422 -4342 332186 -4106
rect 332422 -4342 368186 -4106
rect 368422 -4342 404186 -4106
rect 404422 -4342 440186 -4106
rect 440422 -4342 476186 -4106
rect 476422 -4342 512186 -4106
rect 512422 -4342 548186 -4106
rect 548422 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 8186 -4426
rect 8422 -4662 44186 -4426
rect 44422 -4662 80186 -4426
rect 80422 -4662 116186 -4426
rect 116422 -4662 152186 -4426
rect 152422 -4662 188186 -4426
rect 188422 -4662 224186 -4426
rect 224422 -4662 260186 -4426
rect 260422 -4662 296186 -4426
rect 296422 -4662 332186 -4426
rect 332422 -4662 368186 -4426
rect 368422 -4662 404186 -4426
rect 404422 -4662 440186 -4426
rect 440422 -4662 476186 -4426
rect 476422 -4662 512186 -4426
rect 512422 -4662 548186 -4426
rect 548422 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 152004 -4686 152604 -4684
rect 188004 -4686 188604 -4684
rect 224004 -4686 224604 -4684
rect 260004 -4686 260604 -4684
rect 296004 -4686 296604 -4684
rect 332004 -4686 332604 -4684
rect 368004 -4686 368604 -4684
rect 404004 -4686 404604 -4684
rect 440004 -4686 440604 -4684
rect 476004 -4686 476604 -4684
rect 512004 -4686 512604 -4684
rect 548004 -4686 548604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 134004 -5024 134604 -5022
rect 170004 -5024 170604 -5022
rect 206004 -5024 206604 -5022
rect 242004 -5024 242604 -5022
rect 278004 -5024 278604 -5022
rect 314004 -5024 314604 -5022
rect 350004 -5024 350604 -5022
rect 386004 -5024 386604 -5022
rect 422004 -5024 422604 -5022
rect 458004 -5024 458604 -5022
rect 494004 -5024 494604 -5022
rect 530004 -5024 530604 -5022
rect 566004 -5024 566604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 26186 -5046
rect 26422 -5282 62186 -5046
rect 62422 -5282 98186 -5046
rect 98422 -5282 134186 -5046
rect 134422 -5282 170186 -5046
rect 170422 -5282 206186 -5046
rect 206422 -5282 242186 -5046
rect 242422 -5282 278186 -5046
rect 278422 -5282 314186 -5046
rect 314422 -5282 350186 -5046
rect 350422 -5282 386186 -5046
rect 386422 -5282 422186 -5046
rect 422422 -5282 458186 -5046
rect 458422 -5282 494186 -5046
rect 494422 -5282 530186 -5046
rect 530422 -5282 566186 -5046
rect 566422 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 26186 -5366
rect 26422 -5602 62186 -5366
rect 62422 -5602 98186 -5366
rect 98422 -5602 134186 -5366
rect 134422 -5602 170186 -5366
rect 170422 -5602 206186 -5366
rect 206422 -5602 242186 -5366
rect 242422 -5602 278186 -5366
rect 278422 -5602 314186 -5366
rect 314422 -5602 350186 -5366
rect 350422 -5602 386186 -5366
rect 386422 -5602 422186 -5366
rect 422422 -5602 458186 -5366
rect 458422 -5602 494186 -5366
rect 494422 -5602 530186 -5366
rect 530422 -5602 566186 -5366
rect 566422 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 134004 -5626 134604 -5624
rect 170004 -5626 170604 -5624
rect 206004 -5626 206604 -5624
rect 242004 -5626 242604 -5624
rect 278004 -5626 278604 -5624
rect 314004 -5626 314604 -5624
rect 350004 -5626 350604 -5624
rect 386004 -5626 386604 -5624
rect 422004 -5626 422604 -5624
rect 458004 -5626 458604 -5624
rect 494004 -5626 494604 -5624
rect 530004 -5626 530604 -5624
rect 566004 -5626 566604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 155604 -5964 156204 -5962
rect 191604 -5964 192204 -5962
rect 227604 -5964 228204 -5962
rect 263604 -5964 264204 -5962
rect 299604 -5964 300204 -5962
rect 335604 -5964 336204 -5962
rect 371604 -5964 372204 -5962
rect 407604 -5964 408204 -5962
rect 443604 -5964 444204 -5962
rect 479604 -5964 480204 -5962
rect 515604 -5964 516204 -5962
rect 551604 -5964 552204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 11786 -5986
rect 12022 -6222 47786 -5986
rect 48022 -6222 83786 -5986
rect 84022 -6222 119786 -5986
rect 120022 -6222 155786 -5986
rect 156022 -6222 191786 -5986
rect 192022 -6222 227786 -5986
rect 228022 -6222 263786 -5986
rect 264022 -6222 299786 -5986
rect 300022 -6222 335786 -5986
rect 336022 -6222 371786 -5986
rect 372022 -6222 407786 -5986
rect 408022 -6222 443786 -5986
rect 444022 -6222 479786 -5986
rect 480022 -6222 515786 -5986
rect 516022 -6222 551786 -5986
rect 552022 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 11786 -6306
rect 12022 -6542 47786 -6306
rect 48022 -6542 83786 -6306
rect 84022 -6542 119786 -6306
rect 120022 -6542 155786 -6306
rect 156022 -6542 191786 -6306
rect 192022 -6542 227786 -6306
rect 228022 -6542 263786 -6306
rect 264022 -6542 299786 -6306
rect 300022 -6542 335786 -6306
rect 336022 -6542 371786 -6306
rect 372022 -6542 407786 -6306
rect 408022 -6542 443786 -6306
rect 444022 -6542 479786 -6306
rect 480022 -6542 515786 -6306
rect 516022 -6542 551786 -6306
rect 552022 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 155604 -6566 156204 -6564
rect 191604 -6566 192204 -6564
rect 227604 -6566 228204 -6564
rect 263604 -6566 264204 -6564
rect 299604 -6566 300204 -6564
rect 335604 -6566 336204 -6564
rect 371604 -6566 372204 -6564
rect 407604 -6566 408204 -6564
rect 443604 -6566 444204 -6564
rect 479604 -6566 480204 -6564
rect 515604 -6566 516204 -6564
rect 551604 -6566 552204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 137604 -6904 138204 -6902
rect 173604 -6904 174204 -6902
rect 209604 -6904 210204 -6902
rect 245604 -6904 246204 -6902
rect 281604 -6904 282204 -6902
rect 317604 -6904 318204 -6902
rect 353604 -6904 354204 -6902
rect 389604 -6904 390204 -6902
rect 425604 -6904 426204 -6902
rect 461604 -6904 462204 -6902
rect 497604 -6904 498204 -6902
rect 533604 -6904 534204 -6902
rect 569604 -6904 570204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 29786 -6926
rect 30022 -7162 65786 -6926
rect 66022 -7162 101786 -6926
rect 102022 -7162 137786 -6926
rect 138022 -7162 173786 -6926
rect 174022 -7162 209786 -6926
rect 210022 -7162 245786 -6926
rect 246022 -7162 281786 -6926
rect 282022 -7162 317786 -6926
rect 318022 -7162 353786 -6926
rect 354022 -7162 389786 -6926
rect 390022 -7162 425786 -6926
rect 426022 -7162 461786 -6926
rect 462022 -7162 497786 -6926
rect 498022 -7162 533786 -6926
rect 534022 -7162 569786 -6926
rect 570022 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 29786 -7246
rect 30022 -7482 65786 -7246
rect 66022 -7482 101786 -7246
rect 102022 -7482 137786 -7246
rect 138022 -7482 173786 -7246
rect 174022 -7482 209786 -7246
rect 210022 -7482 245786 -7246
rect 246022 -7482 281786 -7246
rect 282022 -7482 317786 -7246
rect 318022 -7482 353786 -7246
rect 354022 -7482 389786 -7246
rect 390022 -7482 425786 -7246
rect 426022 -7482 461786 -7246
rect 462022 -7482 497786 -7246
rect 498022 -7482 533786 -7246
rect 534022 -7482 569786 -7246
rect 570022 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 137604 -7506 138204 -7504
rect 173604 -7506 174204 -7504
rect 209604 -7506 210204 -7504
rect 245604 -7506 246204 -7504
rect 281604 -7506 282204 -7504
rect 317604 -7506 318204 -7504
rect 353604 -7506 354204 -7504
rect 389604 -7506 390204 -7504
rect 425604 -7506 426204 -7504
rect 461604 -7506 462204 -7504
rect 497604 -7506 498204 -7504
rect 533604 -7506 534204 -7504
rect 569604 -7506 570204 -7504
rect 591900 -7506 592500 -7504
use opamp_v1  opamp_v1_6
timestamp 1606921152
transform -1 0 556309 0 -1 213029
box 2069 -10028 26971 3199
use opamp_v1  opamp_v1_5
timestamp 1606921152
transform -1 0 557443 0 -1 403301
box 2069 -10028 26971 3199
use opamp_v1  opamp_v1_4
timestamp 1606921152
transform -1 0 557481 0 -1 588029
box 2069 -10028 26971 3199
use opamp_v1  opamp_v1_3
timestamp 1606921152
transform 0 1 479026 -1 0 677687
box 2069 -10028 26971 3199
use opamp_v1  opamp_v1_2
timestamp 1606921152
transform 0 1 220266 -1 0 678857
box 2069 -10028 26971 3199
use opamp_v1  opamp_v1_1
timestamp 1606921152
transform 1 0 23845 0 1 611502
box 2069 -10028 26971 3199
use opamp_v1  opamp_v1_0
timestamp 1606921152
transform 1 0 23351 0 1 439806
box 2069 -10028 26971 3199
use PLL_  PLL__0
timestamp 1607692587
transform 1 0 12492 0 1 15176
box -4474 -3468 12028 4060
<< labels >>
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal4 s 576804 703520 577404 705800 6 vccd1
port 636 nsew default input
rlabel metal4 s 540804 703520 541404 705800 6 vccd1
port 637 nsew default input
rlabel metal4 s 504804 703520 505404 705800 6 vccd1
port 638 nsew default input
rlabel metal4 s 468804 703520 469404 705800 6 vccd1
port 639 nsew default input
rlabel metal4 s 432804 703520 433404 705800 6 vccd1
port 640 nsew default input
rlabel metal4 s 396804 703520 397404 705800 6 vccd1
port 641 nsew default input
rlabel metal4 s 360804 703520 361404 705800 6 vccd1
port 642 nsew default input
rlabel metal4 s 324804 703520 325404 705800 6 vccd1
port 643 nsew default input
rlabel metal4 s 288804 703520 289404 705800 6 vccd1
port 644 nsew default input
rlabel metal4 s 252804 703520 253404 705800 6 vccd1
port 645 nsew default input
rlabel metal4 s 216804 703520 217404 705800 6 vccd1
port 646 nsew default input
rlabel metal4 s 180804 703520 181404 705800 6 vccd1
port 647 nsew default input
rlabel metal4 s 144804 703520 145404 705800 6 vccd1
port 648 nsew default input
rlabel metal4 s 108804 703520 109404 705800 6 vccd1
port 649 nsew default input
rlabel metal4 s 72804 703520 73404 705800 6 vccd1
port 650 nsew default input
rlabel metal4 s 36804 703520 37404 705800 6 vccd1
port 651 nsew default input
rlabel metal4 s 804 703520 1404 705800 6 vccd1
port 652 nsew default input
rlabel metal4 s 585320 -924 585920 704860 6 vccd1
port 653 nsew default input
rlabel metal4 s -1996 -924 -1396 704860 4 vccd1
port 654 nsew default input
rlabel metal4 s 576804 -1864 577404 480 8 vccd1
port 655 nsew default input
rlabel metal4 s 540804 -1864 541404 480 8 vccd1
port 656 nsew default input
rlabel metal4 s 504804 -1864 505404 480 8 vccd1
port 657 nsew default input
rlabel metal4 s 468804 -1864 469404 480 8 vccd1
port 658 nsew default input
rlabel metal4 s 432804 -1864 433404 480 8 vccd1
port 659 nsew default input
rlabel metal4 s 396804 -1864 397404 480 8 vccd1
port 660 nsew default input
rlabel metal4 s 360804 -1864 361404 480 8 vccd1
port 661 nsew default input
rlabel metal4 s 324804 -1864 325404 480 8 vccd1
port 662 nsew default input
rlabel metal4 s 288804 -1864 289404 480 8 vccd1
port 663 nsew default input
rlabel metal4 s 252804 -1864 253404 480 8 vccd1
port 664 nsew default input
rlabel metal4 s 216804 -1864 217404 480 8 vccd1
port 665 nsew default input
rlabel metal4 s 180804 -1864 181404 480 8 vccd1
port 666 nsew default input
rlabel metal4 s 144804 -1864 145404 480 8 vccd1
port 667 nsew default input
rlabel metal4 s 108804 -1864 109404 480 8 vccd1
port 668 nsew default input
rlabel metal4 s 72804 -1864 73404 480 8 vccd1
port 669 nsew default input
rlabel metal4 s 36804 -1864 37404 480 8 vccd1
port 670 nsew default input
rlabel metal4 s 804 -1864 1404 480 8 vccd1
port 671 nsew default input
rlabel metal5 s -1996 704260 585920 704860 6 vccd1
port 672 nsew default input
rlabel metal5 s 583520 685876 586860 686476 6 vccd1
port 673 nsew default input
rlabel metal5 s -2936 685876 480 686476 4 vccd1
port 674 nsew default input
rlabel metal5 s 583520 649876 586860 650476 6 vccd1
port 675 nsew default input
rlabel metal5 s -2936 649876 480 650476 4 vccd1
port 676 nsew default input
rlabel metal5 s 583520 613876 586860 614476 6 vccd1
port 677 nsew default input
rlabel metal5 s -2936 613876 480 614476 4 vccd1
port 678 nsew default input
rlabel metal5 s 583520 577876 586860 578476 6 vccd1
port 679 nsew default input
rlabel metal5 s -2936 577876 480 578476 4 vccd1
port 680 nsew default input
rlabel metal5 s 583520 541876 586860 542476 6 vccd1
port 681 nsew default input
rlabel metal5 s -2936 541876 480 542476 4 vccd1
port 682 nsew default input
rlabel metal5 s 583520 505876 586860 506476 6 vccd1
port 683 nsew default input
rlabel metal5 s -2936 505876 480 506476 4 vccd1
port 684 nsew default input
rlabel metal5 s 583520 469876 586860 470476 6 vccd1
port 685 nsew default input
rlabel metal5 s -2936 469876 480 470476 4 vccd1
port 686 nsew default input
rlabel metal5 s 583520 433876 586860 434476 6 vccd1
port 687 nsew default input
rlabel metal5 s -2936 433876 480 434476 4 vccd1
port 688 nsew default input
rlabel metal5 s 583520 397876 586860 398476 6 vccd1
port 689 nsew default input
rlabel metal5 s -2936 397876 480 398476 4 vccd1
port 690 nsew default input
rlabel metal5 s 583520 361876 586860 362476 6 vccd1
port 691 nsew default input
rlabel metal5 s -2936 361876 480 362476 4 vccd1
port 692 nsew default input
rlabel metal5 s 583520 325876 586860 326476 6 vccd1
port 693 nsew default input
rlabel metal5 s -2936 325876 480 326476 4 vccd1
port 694 nsew default input
rlabel metal5 s 583520 289876 586860 290476 6 vccd1
port 695 nsew default input
rlabel metal5 s -2936 289876 480 290476 4 vccd1
port 696 nsew default input
rlabel metal5 s 583520 253876 586860 254476 6 vccd1
port 697 nsew default input
rlabel metal5 s -2936 253876 480 254476 4 vccd1
port 698 nsew default input
rlabel metal5 s 583520 217876 586860 218476 6 vccd1
port 699 nsew default input
rlabel metal5 s -2936 217876 480 218476 4 vccd1
port 700 nsew default input
rlabel metal5 s 583520 181876 586860 182476 6 vccd1
port 701 nsew default input
rlabel metal5 s -2936 181876 480 182476 4 vccd1
port 702 nsew default input
rlabel metal5 s 583520 145876 586860 146476 6 vccd1
port 703 nsew default input
rlabel metal5 s -2936 145876 480 146476 4 vccd1
port 704 nsew default input
rlabel metal5 s 583520 109876 586860 110476 6 vccd1
port 705 nsew default input
rlabel metal5 s -2936 109876 480 110476 4 vccd1
port 706 nsew default input
rlabel metal5 s 583520 73876 586860 74476 6 vccd1
port 707 nsew default input
rlabel metal5 s -2936 73876 480 74476 4 vccd1
port 708 nsew default input
rlabel metal5 s 583520 37876 586860 38476 6 vccd1
port 709 nsew default input
rlabel metal5 s -2936 37876 480 38476 4 vccd1
port 710 nsew default input
rlabel metal5 s 583520 1876 586860 2476 6 vccd1
port 711 nsew default input
rlabel metal5 s -2936 1876 480 2476 4 vccd1
port 712 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 713 nsew default input
rlabel metal4 s 586260 -1864 586860 705800 6 vssd1
port 714 nsew default input
rlabel metal4 s 558804 703520 559404 705800 6 vssd1
port 715 nsew default input
rlabel metal4 s 522804 703520 523404 705800 6 vssd1
port 716 nsew default input
rlabel metal4 s 486804 703520 487404 705800 6 vssd1
port 717 nsew default input
rlabel metal4 s 450804 703520 451404 705800 6 vssd1
port 718 nsew default input
rlabel metal4 s 414804 703520 415404 705800 6 vssd1
port 719 nsew default input
rlabel metal4 s 378804 703520 379404 705800 6 vssd1
port 720 nsew default input
rlabel metal4 s 342804 703520 343404 705800 6 vssd1
port 721 nsew default input
rlabel metal4 s 306804 703520 307404 705800 6 vssd1
port 722 nsew default input
rlabel metal4 s 270804 703520 271404 705800 6 vssd1
port 723 nsew default input
rlabel metal4 s 234804 703520 235404 705800 6 vssd1
port 724 nsew default input
rlabel metal4 s 198804 703520 199404 705800 6 vssd1
port 725 nsew default input
rlabel metal4 s 162804 703520 163404 705800 6 vssd1
port 726 nsew default input
rlabel metal4 s 126804 703520 127404 705800 6 vssd1
port 727 nsew default input
rlabel metal4 s 90804 703520 91404 705800 6 vssd1
port 728 nsew default input
rlabel metal4 s 54804 703520 55404 705800 6 vssd1
port 729 nsew default input
rlabel metal4 s 18804 703520 19404 705800 6 vssd1
port 730 nsew default input
rlabel metal4 s -2936 -1864 -2336 705800 4 vssd1
port 731 nsew default input
rlabel metal4 s 558804 -1864 559404 480 8 vssd1
port 732 nsew default input
rlabel metal4 s 522804 -1864 523404 480 8 vssd1
port 733 nsew default input
rlabel metal4 s 486804 -1864 487404 480 8 vssd1
port 734 nsew default input
rlabel metal4 s 450804 -1864 451404 480 8 vssd1
port 735 nsew default input
rlabel metal4 s 414804 -1864 415404 480 8 vssd1
port 736 nsew default input
rlabel metal4 s 378804 -1864 379404 480 8 vssd1
port 737 nsew default input
rlabel metal4 s 342804 -1864 343404 480 8 vssd1
port 738 nsew default input
rlabel metal4 s 306804 -1864 307404 480 8 vssd1
port 739 nsew default input
rlabel metal4 s 270804 -1864 271404 480 8 vssd1
port 740 nsew default input
rlabel metal4 s 234804 -1864 235404 480 8 vssd1
port 741 nsew default input
rlabel metal4 s 198804 -1864 199404 480 8 vssd1
port 742 nsew default input
rlabel metal4 s 162804 -1864 163404 480 8 vssd1
port 743 nsew default input
rlabel metal4 s 126804 -1864 127404 480 8 vssd1
port 744 nsew default input
rlabel metal4 s 90804 -1864 91404 480 8 vssd1
port 745 nsew default input
rlabel metal4 s 54804 -1864 55404 480 8 vssd1
port 746 nsew default input
rlabel metal4 s 18804 -1864 19404 480 8 vssd1
port 747 nsew default input
rlabel metal5 s -2936 705200 586860 705800 6 vssd1
port 748 nsew default input
rlabel metal5 s 583520 667876 586860 668476 6 vssd1
port 749 nsew default input
rlabel metal5 s -2936 667876 480 668476 4 vssd1
port 750 nsew default input
rlabel metal5 s 583520 631876 586860 632476 6 vssd1
port 751 nsew default input
rlabel metal5 s -2936 631876 480 632476 4 vssd1
port 752 nsew default input
rlabel metal5 s 583520 595876 586860 596476 6 vssd1
port 753 nsew default input
rlabel metal5 s -2936 595876 480 596476 4 vssd1
port 754 nsew default input
rlabel metal5 s 583520 559876 586860 560476 6 vssd1
port 755 nsew default input
rlabel metal5 s -2936 559876 480 560476 4 vssd1
port 756 nsew default input
rlabel metal5 s 583520 523876 586860 524476 6 vssd1
port 757 nsew default input
rlabel metal5 s -2936 523876 480 524476 4 vssd1
port 758 nsew default input
rlabel metal5 s 583520 487876 586860 488476 6 vssd1
port 759 nsew default input
rlabel metal5 s -2936 487876 480 488476 4 vssd1
port 760 nsew default input
rlabel metal5 s 583520 451876 586860 452476 6 vssd1
port 761 nsew default input
rlabel metal5 s -2936 451876 480 452476 4 vssd1
port 762 nsew default input
rlabel metal5 s 583520 415876 586860 416476 6 vssd1
port 763 nsew default input
rlabel metal5 s -2936 415876 480 416476 4 vssd1
port 764 nsew default input
rlabel metal5 s 583520 379876 586860 380476 6 vssd1
port 765 nsew default input
rlabel metal5 s -2936 379876 480 380476 4 vssd1
port 766 nsew default input
rlabel metal5 s 583520 343876 586860 344476 6 vssd1
port 767 nsew default input
rlabel metal5 s -2936 343876 480 344476 4 vssd1
port 768 nsew default input
rlabel metal5 s 583520 307876 586860 308476 6 vssd1
port 769 nsew default input
rlabel metal5 s -2936 307876 480 308476 4 vssd1
port 770 nsew default input
rlabel metal5 s 583520 271876 586860 272476 6 vssd1
port 771 nsew default input
rlabel metal5 s -2936 271876 480 272476 4 vssd1
port 772 nsew default input
rlabel metal5 s 583520 235876 586860 236476 6 vssd1
port 773 nsew default input
rlabel metal5 s -2936 235876 480 236476 4 vssd1
port 774 nsew default input
rlabel metal5 s 583520 199876 586860 200476 6 vssd1
port 775 nsew default input
rlabel metal5 s -2936 199876 480 200476 4 vssd1
port 776 nsew default input
rlabel metal5 s 583520 163876 586860 164476 6 vssd1
port 777 nsew default input
rlabel metal5 s -2936 163876 480 164476 4 vssd1
port 778 nsew default input
rlabel metal5 s 583520 127876 586860 128476 6 vssd1
port 779 nsew default input
rlabel metal5 s -2936 127876 480 128476 4 vssd1
port 780 nsew default input
rlabel metal5 s 583520 91876 586860 92476 6 vssd1
port 781 nsew default input
rlabel metal5 s -2936 91876 480 92476 4 vssd1
port 782 nsew default input
rlabel metal5 s 583520 55876 586860 56476 6 vssd1
port 783 nsew default input
rlabel metal5 s -2936 55876 480 56476 4 vssd1
port 784 nsew default input
rlabel metal5 s 583520 19876 586860 20476 6 vssd1
port 785 nsew default input
rlabel metal5 s -2936 19876 480 20476 4 vssd1
port 786 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 787 nsew default input
rlabel metal4 s 580404 703520 581004 707680 6 vccd2
port 788 nsew default input
rlabel metal4 s 544404 703520 545004 707680 6 vccd2
port 789 nsew default input
rlabel metal4 s 508404 703520 509004 707680 6 vccd2
port 790 nsew default input
rlabel metal4 s 472404 703520 473004 707680 6 vccd2
port 791 nsew default input
rlabel metal4 s 436404 703520 437004 707680 6 vccd2
port 792 nsew default input
rlabel metal4 s 400404 703520 401004 707680 6 vccd2
port 793 nsew default input
rlabel metal4 s 364404 703520 365004 707680 6 vccd2
port 794 nsew default input
rlabel metal4 s 328404 703520 329004 707680 6 vccd2
port 795 nsew default input
rlabel metal4 s 292404 703520 293004 707680 6 vccd2
port 796 nsew default input
rlabel metal4 s 256404 703520 257004 707680 6 vccd2
port 797 nsew default input
rlabel metal4 s 220404 703520 221004 707680 6 vccd2
port 798 nsew default input
rlabel metal4 s 184404 703520 185004 707680 6 vccd2
port 799 nsew default input
rlabel metal4 s 148404 703520 149004 707680 6 vccd2
port 800 nsew default input
rlabel metal4 s 112404 703520 113004 707680 6 vccd2
port 801 nsew default input
rlabel metal4 s 76404 703520 77004 707680 6 vccd2
port 802 nsew default input
rlabel metal4 s 40404 703520 41004 707680 6 vccd2
port 803 nsew default input
rlabel metal4 s 4404 703520 5004 707680 6 vccd2
port 804 nsew default input
rlabel metal4 s 587200 -2804 587800 706740 6 vccd2
port 805 nsew default input
rlabel metal4 s -3876 -2804 -3276 706740 4 vccd2
port 806 nsew default input
rlabel metal4 s 580404 -3744 581004 480 8 vccd2
port 807 nsew default input
rlabel metal4 s 544404 -3744 545004 480 8 vccd2
port 808 nsew default input
rlabel metal4 s 508404 -3744 509004 480 8 vccd2
port 809 nsew default input
rlabel metal4 s 472404 -3744 473004 480 8 vccd2
port 810 nsew default input
rlabel metal4 s 436404 -3744 437004 480 8 vccd2
port 811 nsew default input
rlabel metal4 s 400404 -3744 401004 480 8 vccd2
port 812 nsew default input
rlabel metal4 s 364404 -3744 365004 480 8 vccd2
port 813 nsew default input
rlabel metal4 s 328404 -3744 329004 480 8 vccd2
port 814 nsew default input
rlabel metal4 s 292404 -3744 293004 480 8 vccd2
port 815 nsew default input
rlabel metal4 s 256404 -3744 257004 480 8 vccd2
port 816 nsew default input
rlabel metal4 s 220404 -3744 221004 480 8 vccd2
port 817 nsew default input
rlabel metal4 s 184404 -3744 185004 480 8 vccd2
port 818 nsew default input
rlabel metal4 s 148404 -3744 149004 480 8 vccd2
port 819 nsew default input
rlabel metal4 s 112404 -3744 113004 480 8 vccd2
port 820 nsew default input
rlabel metal4 s 76404 -3744 77004 480 8 vccd2
port 821 nsew default input
rlabel metal4 s 40404 -3744 41004 480 8 vccd2
port 822 nsew default input
rlabel metal4 s 4404 -3744 5004 480 8 vccd2
port 823 nsew default input
rlabel metal5 s -3876 706140 587800 706740 6 vccd2
port 824 nsew default input
rlabel metal5 s 583520 689476 588740 690076 6 vccd2
port 825 nsew default input
rlabel metal5 s -4816 689476 480 690076 4 vccd2
port 826 nsew default input
rlabel metal5 s 583520 653476 588740 654076 6 vccd2
port 827 nsew default input
rlabel metal5 s -4816 653476 480 654076 4 vccd2
port 828 nsew default input
rlabel metal5 s 583520 617476 588740 618076 6 vccd2
port 829 nsew default input
rlabel metal5 s -4816 617476 480 618076 4 vccd2
port 830 nsew default input
rlabel metal5 s 583520 581476 588740 582076 6 vccd2
port 831 nsew default input
rlabel metal5 s -4816 581476 480 582076 4 vccd2
port 832 nsew default input
rlabel metal5 s 583520 545476 588740 546076 6 vccd2
port 833 nsew default input
rlabel metal5 s -4816 545476 480 546076 4 vccd2
port 834 nsew default input
rlabel metal5 s 583520 509476 588740 510076 6 vccd2
port 835 nsew default input
rlabel metal5 s -4816 509476 480 510076 4 vccd2
port 836 nsew default input
rlabel metal5 s 583520 473476 588740 474076 6 vccd2
port 837 nsew default input
rlabel metal5 s -4816 473476 480 474076 4 vccd2
port 838 nsew default input
rlabel metal5 s 583520 437476 588740 438076 6 vccd2
port 839 nsew default input
rlabel metal5 s -4816 437476 480 438076 4 vccd2
port 840 nsew default input
rlabel metal5 s 583520 401476 588740 402076 6 vccd2
port 841 nsew default input
rlabel metal5 s -4816 401476 480 402076 4 vccd2
port 842 nsew default input
rlabel metal5 s 583520 365476 588740 366076 6 vccd2
port 843 nsew default input
rlabel metal5 s -4816 365476 480 366076 4 vccd2
port 844 nsew default input
rlabel metal5 s 583520 329476 588740 330076 6 vccd2
port 845 nsew default input
rlabel metal5 s -4816 329476 480 330076 4 vccd2
port 846 nsew default input
rlabel metal5 s 583520 293476 588740 294076 6 vccd2
port 847 nsew default input
rlabel metal5 s -4816 293476 480 294076 4 vccd2
port 848 nsew default input
rlabel metal5 s 583520 257476 588740 258076 6 vccd2
port 849 nsew default input
rlabel metal5 s -4816 257476 480 258076 4 vccd2
port 850 nsew default input
rlabel metal5 s 583520 221476 588740 222076 6 vccd2
port 851 nsew default input
rlabel metal5 s -4816 221476 480 222076 4 vccd2
port 852 nsew default input
rlabel metal5 s 583520 185476 588740 186076 6 vccd2
port 853 nsew default input
rlabel metal5 s -4816 185476 480 186076 4 vccd2
port 854 nsew default input
rlabel metal5 s 583520 149476 588740 150076 6 vccd2
port 855 nsew default input
rlabel metal5 s -4816 149476 480 150076 4 vccd2
port 856 nsew default input
rlabel metal5 s 583520 113476 588740 114076 6 vccd2
port 857 nsew default input
rlabel metal5 s -4816 113476 480 114076 4 vccd2
port 858 nsew default input
rlabel metal5 s 583520 77476 588740 78076 6 vccd2
port 859 nsew default input
rlabel metal5 s -4816 77476 480 78076 4 vccd2
port 860 nsew default input
rlabel metal5 s 583520 41476 588740 42076 6 vccd2
port 861 nsew default input
rlabel metal5 s -4816 41476 480 42076 4 vccd2
port 862 nsew default input
rlabel metal5 s 583520 5476 588740 6076 6 vccd2
port 863 nsew default input
rlabel metal5 s -4816 5476 480 6076 4 vccd2
port 864 nsew default input
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 865 nsew default input
rlabel metal4 s 588140 -3744 588740 707680 6 vssd2
port 866 nsew default input
rlabel metal4 s 562404 703520 563004 707680 6 vssd2
port 867 nsew default input
rlabel metal4 s 526404 703520 527004 707680 6 vssd2
port 868 nsew default input
rlabel metal4 s 490404 703520 491004 707680 6 vssd2
port 869 nsew default input
rlabel metal4 s 454404 703520 455004 707680 6 vssd2
port 870 nsew default input
rlabel metal4 s 418404 703520 419004 707680 6 vssd2
port 871 nsew default input
rlabel metal4 s 382404 703520 383004 707680 6 vssd2
port 872 nsew default input
rlabel metal4 s 346404 703520 347004 707680 6 vssd2
port 873 nsew default input
rlabel metal4 s 310404 703520 311004 707680 6 vssd2
port 874 nsew default input
rlabel metal4 s 274404 703520 275004 707680 6 vssd2
port 875 nsew default input
rlabel metal4 s 238404 703520 239004 707680 6 vssd2
port 876 nsew default input
rlabel metal4 s 202404 703520 203004 707680 6 vssd2
port 877 nsew default input
rlabel metal4 s 166404 703520 167004 707680 6 vssd2
port 878 nsew default input
rlabel metal4 s 130404 703520 131004 707680 6 vssd2
port 879 nsew default input
rlabel metal4 s 94404 703520 95004 707680 6 vssd2
port 880 nsew default input
rlabel metal4 s 58404 703520 59004 707680 6 vssd2
port 881 nsew default input
rlabel metal4 s 22404 703520 23004 707680 6 vssd2
port 882 nsew default input
rlabel metal4 s -4816 -3744 -4216 707680 4 vssd2
port 883 nsew default input
rlabel metal4 s 562404 -3744 563004 480 8 vssd2
port 884 nsew default input
rlabel metal4 s 526404 -3744 527004 480 8 vssd2
port 885 nsew default input
rlabel metal4 s 490404 -3744 491004 480 8 vssd2
port 886 nsew default input
rlabel metal4 s 454404 -3744 455004 480 8 vssd2
port 887 nsew default input
rlabel metal4 s 418404 -3744 419004 480 8 vssd2
port 888 nsew default input
rlabel metal4 s 382404 -3744 383004 480 8 vssd2
port 889 nsew default input
rlabel metal4 s 346404 -3744 347004 480 8 vssd2
port 890 nsew default input
rlabel metal4 s 310404 -3744 311004 480 8 vssd2
port 891 nsew default input
rlabel metal4 s 274404 -3744 275004 480 8 vssd2
port 892 nsew default input
rlabel metal4 s 238404 -3744 239004 480 8 vssd2
port 893 nsew default input
rlabel metal4 s 202404 -3744 203004 480 8 vssd2
port 894 nsew default input
rlabel metal4 s 166404 -3744 167004 480 8 vssd2
port 895 nsew default input
rlabel metal4 s 130404 -3744 131004 480 8 vssd2
port 896 nsew default input
rlabel metal4 s 94404 -3744 95004 480 8 vssd2
port 897 nsew default input
rlabel metal4 s 58404 -3744 59004 480 8 vssd2
port 898 nsew default input
rlabel metal4 s 22404 -3744 23004 480 8 vssd2
port 899 nsew default input
rlabel metal5 s -4816 707080 588740 707680 6 vssd2
port 900 nsew default input
rlabel metal5 s 583520 671476 588740 672076 6 vssd2
port 901 nsew default input
rlabel metal5 s -4816 671476 480 672076 4 vssd2
port 902 nsew default input
rlabel metal5 s 583520 635476 588740 636076 6 vssd2
port 903 nsew default input
rlabel metal5 s -4816 635476 480 636076 4 vssd2
port 904 nsew default input
rlabel metal5 s 583520 599476 588740 600076 6 vssd2
port 905 nsew default input
rlabel metal5 s -4816 599476 480 600076 4 vssd2
port 906 nsew default input
rlabel metal5 s 583520 563476 588740 564076 6 vssd2
port 907 nsew default input
rlabel metal5 s -4816 563476 480 564076 4 vssd2
port 908 nsew default input
rlabel metal5 s 583520 527476 588740 528076 6 vssd2
port 909 nsew default input
rlabel metal5 s -4816 527476 480 528076 4 vssd2
port 910 nsew default input
rlabel metal5 s 583520 491476 588740 492076 6 vssd2
port 911 nsew default input
rlabel metal5 s -4816 491476 480 492076 4 vssd2
port 912 nsew default input
rlabel metal5 s 583520 455476 588740 456076 6 vssd2
port 913 nsew default input
rlabel metal5 s -4816 455476 480 456076 4 vssd2
port 914 nsew default input
rlabel metal5 s 583520 419476 588740 420076 6 vssd2
port 915 nsew default input
rlabel metal5 s -4816 419476 480 420076 4 vssd2
port 916 nsew default input
rlabel metal5 s 583520 383476 588740 384076 6 vssd2
port 917 nsew default input
rlabel metal5 s -4816 383476 480 384076 4 vssd2
port 918 nsew default input
rlabel metal5 s 583520 347476 588740 348076 6 vssd2
port 919 nsew default input
rlabel metal5 s -4816 347476 480 348076 4 vssd2
port 920 nsew default input
rlabel metal5 s 583520 311476 588740 312076 6 vssd2
port 921 nsew default input
rlabel metal5 s -4816 311476 480 312076 4 vssd2
port 922 nsew default input
rlabel metal5 s 583520 275476 588740 276076 6 vssd2
port 923 nsew default input
rlabel metal5 s -4816 275476 480 276076 4 vssd2
port 924 nsew default input
rlabel metal5 s 583520 239476 588740 240076 6 vssd2
port 925 nsew default input
rlabel metal5 s -4816 239476 480 240076 4 vssd2
port 926 nsew default input
rlabel metal5 s 583520 203476 588740 204076 6 vssd2
port 927 nsew default input
rlabel metal5 s -4816 203476 480 204076 4 vssd2
port 928 nsew default input
rlabel metal5 s 583520 167476 588740 168076 6 vssd2
port 929 nsew default input
rlabel metal5 s -4816 167476 480 168076 4 vssd2
port 930 nsew default input
rlabel metal5 s 583520 131476 588740 132076 6 vssd2
port 931 nsew default input
rlabel metal5 s -4816 131476 480 132076 4 vssd2
port 932 nsew default input
rlabel metal5 s 583520 95476 588740 96076 6 vssd2
port 933 nsew default input
rlabel metal5 s -4816 95476 480 96076 4 vssd2
port 934 nsew default input
rlabel metal5 s 583520 59476 588740 60076 6 vssd2
port 935 nsew default input
rlabel metal5 s -4816 59476 480 60076 4 vssd2
port 936 nsew default input
rlabel metal5 s 583520 23476 588740 24076 6 vssd2
port 937 nsew default input
rlabel metal5 s -4816 23476 480 24076 4 vssd2
port 938 nsew default input
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 939 nsew default input
rlabel metal4 s 548004 703520 548604 709560 6 vdda1
port 940 nsew default input
rlabel metal4 s 512004 703520 512604 709560 6 vdda1
port 941 nsew default input
rlabel metal4 s 476004 703520 476604 709560 6 vdda1
port 942 nsew default input
rlabel metal4 s 440004 703520 440604 709560 6 vdda1
port 943 nsew default input
rlabel metal4 s 404004 703520 404604 709560 6 vdda1
port 944 nsew default input
rlabel metal4 s 368004 703520 368604 709560 6 vdda1
port 945 nsew default input
rlabel metal4 s 332004 703520 332604 709560 6 vdda1
port 946 nsew default input
rlabel metal4 s 296004 703520 296604 709560 6 vdda1
port 947 nsew default input
rlabel metal4 s 260004 703520 260604 709560 6 vdda1
port 948 nsew default input
rlabel metal4 s 224004 703520 224604 709560 6 vdda1
port 949 nsew default input
rlabel metal4 s 188004 703520 188604 709560 6 vdda1
port 950 nsew default input
rlabel metal4 s 152004 703520 152604 709560 6 vdda1
port 951 nsew default input
rlabel metal4 s 116004 703520 116604 709560 6 vdda1
port 952 nsew default input
rlabel metal4 s 80004 703520 80604 709560 6 vdda1
port 953 nsew default input
rlabel metal4 s 44004 703520 44604 709560 6 vdda1
port 954 nsew default input
rlabel metal4 s 8004 703520 8604 709560 6 vdda1
port 955 nsew default input
rlabel metal4 s 589080 -4684 589680 708620 6 vdda1
port 956 nsew default input
rlabel metal4 s -5756 -4684 -5156 708620 4 vdda1
port 957 nsew default input
rlabel metal4 s 548004 -5624 548604 480 8 vdda1
port 958 nsew default input
rlabel metal4 s 512004 -5624 512604 480 8 vdda1
port 959 nsew default input
rlabel metal4 s 476004 -5624 476604 480 8 vdda1
port 960 nsew default input
rlabel metal4 s 440004 -5624 440604 480 8 vdda1
port 961 nsew default input
rlabel metal4 s 404004 -5624 404604 480 8 vdda1
port 962 nsew default input
rlabel metal4 s 368004 -5624 368604 480 8 vdda1
port 963 nsew default input
rlabel metal4 s 332004 -5624 332604 480 8 vdda1
port 964 nsew default input
rlabel metal4 s 296004 -5624 296604 480 8 vdda1
port 965 nsew default input
rlabel metal4 s 260004 -5624 260604 480 8 vdda1
port 966 nsew default input
rlabel metal4 s 224004 -5624 224604 480 8 vdda1
port 967 nsew default input
rlabel metal4 s 188004 -5624 188604 480 8 vdda1
port 968 nsew default input
rlabel metal4 s 152004 -5624 152604 480 8 vdda1
port 969 nsew default input
rlabel metal4 s 116004 -5624 116604 480 8 vdda1
port 970 nsew default input
rlabel metal4 s 80004 -5624 80604 480 8 vdda1
port 971 nsew default input
rlabel metal4 s 44004 -5624 44604 480 8 vdda1
port 972 nsew default input
rlabel metal4 s 8004 -5624 8604 480 8 vdda1
port 973 nsew default input
rlabel metal5 s -5756 708020 589680 708620 6 vdda1
port 974 nsew default input
rlabel metal5 s 583520 693076 590620 693676 6 vdda1
port 975 nsew default input
rlabel metal5 s -6696 693076 480 693676 4 vdda1
port 976 nsew default input
rlabel metal5 s 583520 657076 590620 657676 6 vdda1
port 977 nsew default input
rlabel metal5 s -6696 657076 480 657676 4 vdda1
port 978 nsew default input
rlabel metal5 s 583520 621076 590620 621676 6 vdda1
port 979 nsew default input
rlabel metal5 s -6696 621076 480 621676 4 vdda1
port 980 nsew default input
rlabel metal5 s 583520 585076 590620 585676 6 vdda1
port 981 nsew default input
rlabel metal5 s -6696 585076 480 585676 4 vdda1
port 982 nsew default input
rlabel metal5 s 583520 549076 590620 549676 6 vdda1
port 983 nsew default input
rlabel metal5 s -6696 549076 480 549676 4 vdda1
port 984 nsew default input
rlabel metal5 s 583520 513076 590620 513676 6 vdda1
port 985 nsew default input
rlabel metal5 s -6696 513076 480 513676 4 vdda1
port 986 nsew default input
rlabel metal5 s 583520 477076 590620 477676 6 vdda1
port 987 nsew default input
rlabel metal5 s -6696 477076 480 477676 4 vdda1
port 988 nsew default input
rlabel metal5 s 583520 441076 590620 441676 6 vdda1
port 989 nsew default input
rlabel metal5 s -6696 441076 480 441676 4 vdda1
port 990 nsew default input
rlabel metal5 s 583520 405076 590620 405676 6 vdda1
port 991 nsew default input
rlabel metal5 s -6696 405076 480 405676 4 vdda1
port 992 nsew default input
rlabel metal5 s 583520 369076 590620 369676 6 vdda1
port 993 nsew default input
rlabel metal5 s -6696 369076 480 369676 4 vdda1
port 994 nsew default input
rlabel metal5 s 583520 333076 590620 333676 6 vdda1
port 995 nsew default input
rlabel metal5 s -6696 333076 480 333676 4 vdda1
port 996 nsew default input
rlabel metal5 s 583520 297076 590620 297676 6 vdda1
port 997 nsew default input
rlabel metal5 s -6696 297076 480 297676 4 vdda1
port 998 nsew default input
rlabel metal5 s 583520 261076 590620 261676 6 vdda1
port 999 nsew default input
rlabel metal5 s -6696 261076 480 261676 4 vdda1
port 1000 nsew default input
rlabel metal5 s 583520 225076 590620 225676 6 vdda1
port 1001 nsew default input
rlabel metal5 s -6696 225076 480 225676 4 vdda1
port 1002 nsew default input
rlabel metal5 s 583520 189076 590620 189676 6 vdda1
port 1003 nsew default input
rlabel metal5 s -6696 189076 480 189676 4 vdda1
port 1004 nsew default input
rlabel metal5 s 583520 153076 590620 153676 6 vdda1
port 1005 nsew default input
rlabel metal5 s -6696 153076 480 153676 4 vdda1
port 1006 nsew default input
rlabel metal5 s 583520 117076 590620 117676 6 vdda1
port 1007 nsew default input
rlabel metal5 s -6696 117076 480 117676 4 vdda1
port 1008 nsew default input
rlabel metal5 s 583520 81076 590620 81676 6 vdda1
port 1009 nsew default input
rlabel metal5 s -6696 81076 480 81676 4 vdda1
port 1010 nsew default input
rlabel metal5 s 583520 45076 590620 45676 6 vdda1
port 1011 nsew default input
rlabel metal5 s -6696 45076 480 45676 4 vdda1
port 1012 nsew default input
rlabel metal5 s 583520 9076 590620 9676 6 vdda1
port 1013 nsew default input
rlabel metal5 s -6696 9076 480 9676 4 vdda1
port 1014 nsew default input
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 1015 nsew default input
rlabel metal4 s 590020 -5624 590620 709560 6 vssa1
port 1016 nsew default input
rlabel metal4 s 566004 703520 566604 709560 6 vssa1
port 1017 nsew default input
rlabel metal4 s 530004 703520 530604 709560 6 vssa1
port 1018 nsew default input
rlabel metal4 s 494004 703520 494604 709560 6 vssa1
port 1019 nsew default input
rlabel metal4 s 458004 703520 458604 709560 6 vssa1
port 1020 nsew default input
rlabel metal4 s 422004 703520 422604 709560 6 vssa1
port 1021 nsew default input
rlabel metal4 s 386004 703520 386604 709560 6 vssa1
port 1022 nsew default input
rlabel metal4 s 350004 703520 350604 709560 6 vssa1
port 1023 nsew default input
rlabel metal4 s 314004 703520 314604 709560 6 vssa1
port 1024 nsew default input
rlabel metal4 s 278004 703520 278604 709560 6 vssa1
port 1025 nsew default input
rlabel metal4 s 242004 703520 242604 709560 6 vssa1
port 1026 nsew default input
rlabel metal4 s 206004 703520 206604 709560 6 vssa1
port 1027 nsew default input
rlabel metal4 s 170004 703520 170604 709560 6 vssa1
port 1028 nsew default input
rlabel metal4 s 134004 703520 134604 709560 6 vssa1
port 1029 nsew default input
rlabel metal4 s 98004 703520 98604 709560 6 vssa1
port 1030 nsew default input
rlabel metal4 s 62004 703520 62604 709560 6 vssa1
port 1031 nsew default input
rlabel metal4 s 26004 703520 26604 709560 6 vssa1
port 1032 nsew default input
rlabel metal4 s -6696 -5624 -6096 709560 4 vssa1
port 1033 nsew default input
rlabel metal4 s 566004 -5624 566604 480 8 vssa1
port 1034 nsew default input
rlabel metal4 s 530004 -5624 530604 480 8 vssa1
port 1035 nsew default input
rlabel metal4 s 494004 -5624 494604 480 8 vssa1
port 1036 nsew default input
rlabel metal4 s 458004 -5624 458604 480 8 vssa1
port 1037 nsew default input
rlabel metal4 s 422004 -5624 422604 480 8 vssa1
port 1038 nsew default input
rlabel metal4 s 386004 -5624 386604 480 8 vssa1
port 1039 nsew default input
rlabel metal4 s 350004 -5624 350604 480 8 vssa1
port 1040 nsew default input
rlabel metal4 s 314004 -5624 314604 480 8 vssa1
port 1041 nsew default input
rlabel metal4 s 278004 -5624 278604 480 8 vssa1
port 1042 nsew default input
rlabel metal4 s 242004 -5624 242604 480 8 vssa1
port 1043 nsew default input
rlabel metal4 s 206004 -5624 206604 480 8 vssa1
port 1044 nsew default input
rlabel metal4 s 170004 -5624 170604 480 8 vssa1
port 1045 nsew default input
rlabel metal4 s 134004 -5624 134604 480 8 vssa1
port 1046 nsew default input
rlabel metal4 s 98004 -5624 98604 480 8 vssa1
port 1047 nsew default input
rlabel metal4 s 62004 -5624 62604 480 8 vssa1
port 1048 nsew default input
rlabel metal4 s 26004 -5624 26604 480 8 vssa1
port 1049 nsew default input
rlabel metal5 s -6696 708960 590620 709560 6 vssa1
port 1050 nsew default input
rlabel metal5 s 583520 675076 590620 675676 6 vssa1
port 1051 nsew default input
rlabel metal5 s -6696 675076 480 675676 4 vssa1
port 1052 nsew default input
rlabel metal5 s 583520 639076 590620 639676 6 vssa1
port 1053 nsew default input
rlabel metal5 s -6696 639076 480 639676 4 vssa1
port 1054 nsew default input
rlabel metal5 s 583520 603076 590620 603676 6 vssa1
port 1055 nsew default input
rlabel metal5 s -6696 603076 480 603676 4 vssa1
port 1056 nsew default input
rlabel metal5 s 583520 567076 590620 567676 6 vssa1
port 1057 nsew default input
rlabel metal5 s -6696 567076 480 567676 4 vssa1
port 1058 nsew default input
rlabel metal5 s 583520 531076 590620 531676 6 vssa1
port 1059 nsew default input
rlabel metal5 s -6696 531076 480 531676 4 vssa1
port 1060 nsew default input
rlabel metal5 s 583520 495076 590620 495676 6 vssa1
port 1061 nsew default input
rlabel metal5 s -6696 495076 480 495676 4 vssa1
port 1062 nsew default input
rlabel metal5 s 583520 459076 590620 459676 6 vssa1
port 1063 nsew default input
rlabel metal5 s -6696 459076 480 459676 4 vssa1
port 1064 nsew default input
rlabel metal5 s 583520 423076 590620 423676 6 vssa1
port 1065 nsew default input
rlabel metal5 s -6696 423076 480 423676 4 vssa1
port 1066 nsew default input
rlabel metal5 s 583520 387076 590620 387676 6 vssa1
port 1067 nsew default input
rlabel metal5 s -6696 387076 480 387676 4 vssa1
port 1068 nsew default input
rlabel metal5 s 583520 351076 590620 351676 6 vssa1
port 1069 nsew default input
rlabel metal5 s -6696 351076 480 351676 4 vssa1
port 1070 nsew default input
rlabel metal5 s 583520 315076 590620 315676 6 vssa1
port 1071 nsew default input
rlabel metal5 s -6696 315076 480 315676 4 vssa1
port 1072 nsew default input
rlabel metal5 s 583520 279076 590620 279676 6 vssa1
port 1073 nsew default input
rlabel metal5 s -6696 279076 480 279676 4 vssa1
port 1074 nsew default input
rlabel metal5 s 583520 243076 590620 243676 6 vssa1
port 1075 nsew default input
rlabel metal5 s -6696 243076 480 243676 4 vssa1
port 1076 nsew default input
rlabel metal5 s 583520 207076 590620 207676 6 vssa1
port 1077 nsew default input
rlabel metal5 s -6696 207076 480 207676 4 vssa1
port 1078 nsew default input
rlabel metal5 s 583520 171076 590620 171676 6 vssa1
port 1079 nsew default input
rlabel metal5 s -6696 171076 480 171676 4 vssa1
port 1080 nsew default input
rlabel metal5 s 583520 135076 590620 135676 6 vssa1
port 1081 nsew default input
rlabel metal5 s -6696 135076 480 135676 4 vssa1
port 1082 nsew default input
rlabel metal5 s 583520 99076 590620 99676 6 vssa1
port 1083 nsew default input
rlabel metal5 s -6696 99076 480 99676 4 vssa1
port 1084 nsew default input
rlabel metal5 s 583520 63076 590620 63676 6 vssa1
port 1085 nsew default input
rlabel metal5 s -6696 63076 480 63676 4 vssa1
port 1086 nsew default input
rlabel metal5 s 583520 27076 590620 27676 6 vssa1
port 1087 nsew default input
rlabel metal5 s -6696 27076 480 27676 4 vssa1
port 1088 nsew default input
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 1089 nsew default input
rlabel metal4 s 551604 703520 552204 711440 6 vdda2
port 1090 nsew default input
rlabel metal4 s 515604 703520 516204 711440 6 vdda2
port 1091 nsew default input
rlabel metal4 s 479604 703520 480204 711440 6 vdda2
port 1092 nsew default input
rlabel metal4 s 443604 703520 444204 711440 6 vdda2
port 1093 nsew default input
rlabel metal4 s 407604 703520 408204 711440 6 vdda2
port 1094 nsew default input
rlabel metal4 s 371604 703520 372204 711440 6 vdda2
port 1095 nsew default input
rlabel metal4 s 335604 703520 336204 711440 6 vdda2
port 1096 nsew default input
rlabel metal4 s 299604 703520 300204 711440 6 vdda2
port 1097 nsew default input
rlabel metal4 s 263604 703520 264204 711440 6 vdda2
port 1098 nsew default input
rlabel metal4 s 227604 703520 228204 711440 6 vdda2
port 1099 nsew default input
rlabel metal4 s 191604 703520 192204 711440 6 vdda2
port 1100 nsew default input
rlabel metal4 s 155604 703520 156204 711440 6 vdda2
port 1101 nsew default input
rlabel metal4 s 119604 703520 120204 711440 6 vdda2
port 1102 nsew default input
rlabel metal4 s 83604 703520 84204 711440 6 vdda2
port 1103 nsew default input
rlabel metal4 s 47604 703520 48204 711440 6 vdda2
port 1104 nsew default input
rlabel metal4 s 11604 703520 12204 711440 6 vdda2
port 1105 nsew default input
rlabel metal4 s 590960 -6564 591560 710500 6 vdda2
port 1106 nsew default input
rlabel metal4 s -7636 -6564 -7036 710500 4 vdda2
port 1107 nsew default input
rlabel metal4 s 551604 -7504 552204 480 8 vdda2
port 1108 nsew default input
rlabel metal4 s 515604 -7504 516204 480 8 vdda2
port 1109 nsew default input
rlabel metal4 s 479604 -7504 480204 480 8 vdda2
port 1110 nsew default input
rlabel metal4 s 443604 -7504 444204 480 8 vdda2
port 1111 nsew default input
rlabel metal4 s 407604 -7504 408204 480 8 vdda2
port 1112 nsew default input
rlabel metal4 s 371604 -7504 372204 480 8 vdda2
port 1113 nsew default input
rlabel metal4 s 335604 -7504 336204 480 8 vdda2
port 1114 nsew default input
rlabel metal4 s 299604 -7504 300204 480 8 vdda2
port 1115 nsew default input
rlabel metal4 s 263604 -7504 264204 480 8 vdda2
port 1116 nsew default input
rlabel metal4 s 227604 -7504 228204 480 8 vdda2
port 1117 nsew default input
rlabel metal4 s 191604 -7504 192204 480 8 vdda2
port 1118 nsew default input
rlabel metal4 s 155604 -7504 156204 480 8 vdda2
port 1119 nsew default input
rlabel metal4 s 119604 -7504 120204 480 8 vdda2
port 1120 nsew default input
rlabel metal4 s 83604 -7504 84204 480 8 vdda2
port 1121 nsew default input
rlabel metal4 s 47604 -7504 48204 480 8 vdda2
port 1122 nsew default input
rlabel metal4 s 11604 -7504 12204 480 8 vdda2
port 1123 nsew default input
rlabel metal5 s -7636 709900 591560 710500 6 vdda2
port 1124 nsew default input
rlabel metal5 s 583520 696676 592500 697276 6 vdda2
port 1125 nsew default input
rlabel metal5 s -8576 696676 480 697276 4 vdda2
port 1126 nsew default input
rlabel metal5 s 583520 660676 592500 661276 6 vdda2
port 1127 nsew default input
rlabel metal5 s -8576 660676 480 661276 4 vdda2
port 1128 nsew default input
rlabel metal5 s 583520 624676 592500 625276 6 vdda2
port 1129 nsew default input
rlabel metal5 s -8576 624676 480 625276 4 vdda2
port 1130 nsew default input
rlabel metal5 s 583520 588676 592500 589276 6 vdda2
port 1131 nsew default input
rlabel metal5 s -8576 588676 480 589276 4 vdda2
port 1132 nsew default input
rlabel metal5 s 583520 552676 592500 553276 6 vdda2
port 1133 nsew default input
rlabel metal5 s -8576 552676 480 553276 4 vdda2
port 1134 nsew default input
rlabel metal5 s 583520 516676 592500 517276 6 vdda2
port 1135 nsew default input
rlabel metal5 s -8576 516676 480 517276 4 vdda2
port 1136 nsew default input
rlabel metal5 s 583520 480676 592500 481276 6 vdda2
port 1137 nsew default input
rlabel metal5 s -8576 480676 480 481276 4 vdda2
port 1138 nsew default input
rlabel metal5 s 583520 444676 592500 445276 6 vdda2
port 1139 nsew default input
rlabel metal5 s -8576 444676 480 445276 4 vdda2
port 1140 nsew default input
rlabel metal5 s 583520 408676 592500 409276 6 vdda2
port 1141 nsew default input
rlabel metal5 s -8576 408676 480 409276 4 vdda2
port 1142 nsew default input
rlabel metal5 s 583520 372676 592500 373276 6 vdda2
port 1143 nsew default input
rlabel metal5 s -8576 372676 480 373276 4 vdda2
port 1144 nsew default input
rlabel metal5 s 583520 336676 592500 337276 6 vdda2
port 1145 nsew default input
rlabel metal5 s -8576 336676 480 337276 4 vdda2
port 1146 nsew default input
rlabel metal5 s 583520 300676 592500 301276 6 vdda2
port 1147 nsew default input
rlabel metal5 s -8576 300676 480 301276 4 vdda2
port 1148 nsew default input
rlabel metal5 s 583520 264676 592500 265276 6 vdda2
port 1149 nsew default input
rlabel metal5 s -8576 264676 480 265276 4 vdda2
port 1150 nsew default input
rlabel metal5 s 583520 228676 592500 229276 6 vdda2
port 1151 nsew default input
rlabel metal5 s -8576 228676 480 229276 4 vdda2
port 1152 nsew default input
rlabel metal5 s 583520 192676 592500 193276 6 vdda2
port 1153 nsew default input
rlabel metal5 s -8576 192676 480 193276 4 vdda2
port 1154 nsew default input
rlabel metal5 s 583520 156676 592500 157276 6 vdda2
port 1155 nsew default input
rlabel metal5 s -8576 156676 480 157276 4 vdda2
port 1156 nsew default input
rlabel metal5 s 583520 120676 592500 121276 6 vdda2
port 1157 nsew default input
rlabel metal5 s -8576 120676 480 121276 4 vdda2
port 1158 nsew default input
rlabel metal5 s 583520 84676 592500 85276 6 vdda2
port 1159 nsew default input
rlabel metal5 s -8576 84676 480 85276 4 vdda2
port 1160 nsew default input
rlabel metal5 s 583520 48676 592500 49276 6 vdda2
port 1161 nsew default input
rlabel metal5 s -8576 48676 480 49276 4 vdda2
port 1162 nsew default input
rlabel metal5 s 583520 12676 592500 13276 6 vdda2
port 1163 nsew default input
rlabel metal5 s -8576 12676 480 13276 4 vdda2
port 1164 nsew default input
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 1165 nsew default input
rlabel metal4 s 591900 -7504 592500 711440 6 vssa2
port 1166 nsew default input
rlabel metal4 s 569604 703520 570204 711440 6 vssa2
port 1167 nsew default input
rlabel metal4 s 533604 703520 534204 711440 6 vssa2
port 1168 nsew default input
rlabel metal4 s 497604 703520 498204 711440 6 vssa2
port 1169 nsew default input
rlabel metal4 s 461604 703520 462204 711440 6 vssa2
port 1170 nsew default input
rlabel metal4 s 425604 703520 426204 711440 6 vssa2
port 1171 nsew default input
rlabel metal4 s 389604 703520 390204 711440 6 vssa2
port 1172 nsew default input
rlabel metal4 s 353604 703520 354204 711440 6 vssa2
port 1173 nsew default input
rlabel metal4 s 317604 703520 318204 711440 6 vssa2
port 1174 nsew default input
rlabel metal4 s 281604 703520 282204 711440 6 vssa2
port 1175 nsew default input
rlabel metal4 s 245604 703520 246204 711440 6 vssa2
port 1176 nsew default input
rlabel metal4 s 209604 703520 210204 711440 6 vssa2
port 1177 nsew default input
rlabel metal4 s 173604 703520 174204 711440 6 vssa2
port 1178 nsew default input
rlabel metal4 s 137604 703520 138204 711440 6 vssa2
port 1179 nsew default input
rlabel metal4 s 101604 703520 102204 711440 6 vssa2
port 1180 nsew default input
rlabel metal4 s 65604 703520 66204 711440 6 vssa2
port 1181 nsew default input
rlabel metal4 s 29604 703520 30204 711440 6 vssa2
port 1182 nsew default input
rlabel metal4 s -8576 -7504 -7976 711440 4 vssa2
port 1183 nsew default input
rlabel metal4 s 569604 -7504 570204 480 8 vssa2
port 1184 nsew default input
rlabel metal4 s 533604 -7504 534204 480 8 vssa2
port 1185 nsew default input
rlabel metal4 s 497604 -7504 498204 480 8 vssa2
port 1186 nsew default input
rlabel metal4 s 461604 -7504 462204 480 8 vssa2
port 1187 nsew default input
rlabel metal4 s 425604 -7504 426204 480 8 vssa2
port 1188 nsew default input
rlabel metal4 s 389604 -7504 390204 480 8 vssa2
port 1189 nsew default input
rlabel metal4 s 353604 -7504 354204 480 8 vssa2
port 1190 nsew default input
rlabel metal4 s 317604 -7504 318204 480 8 vssa2
port 1191 nsew default input
rlabel metal4 s 281604 -7504 282204 480 8 vssa2
port 1192 nsew default input
rlabel metal4 s 245604 -7504 246204 480 8 vssa2
port 1193 nsew default input
rlabel metal4 s 209604 -7504 210204 480 8 vssa2
port 1194 nsew default input
rlabel metal4 s 173604 -7504 174204 480 8 vssa2
port 1195 nsew default input
rlabel metal4 s 137604 -7504 138204 480 8 vssa2
port 1196 nsew default input
rlabel metal4 s 101604 -7504 102204 480 8 vssa2
port 1197 nsew default input
rlabel metal4 s 65604 -7504 66204 480 8 vssa2
port 1198 nsew default input
rlabel metal4 s 29604 -7504 30204 480 8 vssa2
port 1199 nsew default input
rlabel metal5 s -8576 710840 592500 711440 6 vssa2
port 1200 nsew default input
rlabel metal5 s 583520 678676 592500 679276 6 vssa2
port 1201 nsew default input
rlabel metal5 s -8576 678676 480 679276 4 vssa2
port 1202 nsew default input
rlabel metal5 s 583520 642676 592500 643276 6 vssa2
port 1203 nsew default input
rlabel metal5 s -8576 642676 480 643276 4 vssa2
port 1204 nsew default input
rlabel metal5 s 583520 606676 592500 607276 6 vssa2
port 1205 nsew default input
rlabel metal5 s -8576 606676 480 607276 4 vssa2
port 1206 nsew default input
rlabel metal5 s 583520 570676 592500 571276 6 vssa2
port 1207 nsew default input
rlabel metal5 s -8576 570676 480 571276 4 vssa2
port 1208 nsew default input
rlabel metal5 s 583520 534676 592500 535276 6 vssa2
port 1209 nsew default input
rlabel metal5 s -8576 534676 480 535276 4 vssa2
port 1210 nsew default input
rlabel metal5 s 583520 498676 592500 499276 6 vssa2
port 1211 nsew default input
rlabel metal5 s -8576 498676 480 499276 4 vssa2
port 1212 nsew default input
rlabel metal5 s 583520 462676 592500 463276 6 vssa2
port 1213 nsew default input
rlabel metal5 s -8576 462676 480 463276 4 vssa2
port 1214 nsew default input
rlabel metal5 s 583520 426676 592500 427276 6 vssa2
port 1215 nsew default input
rlabel metal5 s -8576 426676 480 427276 4 vssa2
port 1216 nsew default input
rlabel metal5 s 583520 390676 592500 391276 6 vssa2
port 1217 nsew default input
rlabel metal5 s -8576 390676 480 391276 4 vssa2
port 1218 nsew default input
rlabel metal5 s 583520 354676 592500 355276 6 vssa2
port 1219 nsew default input
rlabel metal5 s -8576 354676 480 355276 4 vssa2
port 1220 nsew default input
rlabel metal5 s 583520 318676 592500 319276 6 vssa2
port 1221 nsew default input
rlabel metal5 s -8576 318676 480 319276 4 vssa2
port 1222 nsew default input
rlabel metal5 s 583520 282676 592500 283276 6 vssa2
port 1223 nsew default input
rlabel metal5 s -8576 282676 480 283276 4 vssa2
port 1224 nsew default input
rlabel metal5 s 583520 246676 592500 247276 6 vssa2
port 1225 nsew default input
rlabel metal5 s -8576 246676 480 247276 4 vssa2
port 1226 nsew default input
rlabel metal5 s 583520 210676 592500 211276 6 vssa2
port 1227 nsew default input
rlabel metal5 s -8576 210676 480 211276 4 vssa2
port 1228 nsew default input
rlabel metal5 s 583520 174676 592500 175276 6 vssa2
port 1229 nsew default input
rlabel metal5 s -8576 174676 480 175276 4 vssa2
port 1230 nsew default input
rlabel metal5 s 583520 138676 592500 139276 6 vssa2
port 1231 nsew default input
rlabel metal5 s -8576 138676 480 139276 4 vssa2
port 1232 nsew default input
rlabel metal5 s 583520 102676 592500 103276 6 vssa2
port 1233 nsew default input
rlabel metal5 s -8576 102676 480 103276 4 vssa2
port 1234 nsew default input
rlabel metal5 s 583520 66676 592500 67276 6 vssa2
port 1235 nsew default input
rlabel metal5 s -8576 66676 480 67276 4 vssa2
port 1236 nsew default input
rlabel metal5 s 583520 30676 592500 31276 6 vssa2
port 1237 nsew default input
rlabel metal5 s -8576 30676 480 31276 4 vssa2
port 1238 nsew default input
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 1239 nsew default input
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
