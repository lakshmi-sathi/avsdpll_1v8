magic
tech sky130A
magscale 1 2
timestamp 1607692587
<< locali >>
rect -1296 3182 -1126 3204
rect -1296 3076 -1264 3182
rect -1158 3180 -1126 3182
rect 1858 3184 3396 3196
rect -1158 3152 -178 3180
rect 1858 3152 3398 3184
rect 5458 3152 6596 3204
rect -1158 3118 -56 3152
rect 1734 3118 3548 3152
rect 5354 3118 6716 3152
rect 8516 3118 9170 3164
rect -1158 3076 -178 3118
rect -1296 3050 -178 3076
rect 1858 3080 3398 3118
rect 1858 3064 3396 3080
rect 5458 3064 6596 3118
rect -1296 3048 -1108 3050
rect 9006 2684 9170 3118
rect 11356 3098 11502 3124
rect 11198 3084 11502 3098
rect 11198 3058 11381 3084
rect 11356 3050 11381 3058
rect 11415 3050 11457 3084
rect 11491 3050 11502 3084
rect 11356 3010 11502 3050
rect 9006 2682 9368 2684
rect 9006 2640 9494 2682
rect 9006 2534 9224 2640
rect 9330 2636 9494 2640
rect 9330 2534 9368 2636
rect 9006 2498 9368 2534
rect 9998 1303 10076 1322
rect 9998 1269 10020 1303
rect 10054 1269 10076 1303
rect 9998 1250 10076 1269
rect 10040 1170 10074 1250
rect 3072 1073 3160 1102
rect 3072 1039 3096 1073
rect 3130 1062 3160 1073
rect 8864 1065 9006 1112
rect 3130 1039 3324 1062
rect 3072 1014 3324 1039
rect 8864 1031 8884 1065
rect 8918 1031 8956 1065
rect 8990 1031 9006 1065
rect 8864 982 9006 1031
rect 846 946 952 950
rect 690 912 952 946
rect 846 910 952 912
rect 846 876 883 910
rect 917 876 952 910
rect 846 846 952 876
rect 8874 856 8980 982
rect 7212 750 8980 856
rect 1546 584 1722 586
rect 814 534 1722 584
rect -1992 480 -1662 512
rect 814 498 1594 534
rect -1992 374 -1974 480
rect -1724 398 -1662 480
rect -1724 374 -1110 398
rect -1992 340 -1110 374
rect -1992 338 -1662 340
rect 816 330 894 498
rect 1546 428 1594 498
rect 1700 428 1722 534
rect 1546 402 1722 428
rect 730 296 894 330
rect 8058 -700 8446 750
rect 8784 -700 8828 -698
rect 8058 -930 8828 -700
rect 8606 -962 8828 -930
rect 8606 -1764 8826 -962
rect -384 -1966 -146 -1882
rect 120 -1956 382 -1870
rect 3722 -1958 3952 -1872
rect 4218 -1954 4492 -1868
rect 7840 -1956 8098 -1872
rect 8364 -1984 8826 -1764
<< viali >>
rect -1264 3076 -1158 3182
rect 11381 3050 11415 3084
rect 11457 3050 11491 3084
rect 9224 2534 9330 2640
rect 10020 1269 10054 1303
rect 3096 1039 3130 1073
rect 8884 1031 8918 1065
rect 8956 1031 8990 1065
rect 883 876 917 910
rect -1974 374 -1724 480
rect 1594 428 1700 534
<< metal1 >>
rect -4450 3496 -4336 3568
rect -4450 3400 14 3496
rect 1670 3400 3584 3496
rect 5276 3400 6710 3496
rect 8440 3400 9518 3496
rect -4450 3330 -4336 3400
rect 9272 3237 9416 3252
rect -1322 3189 -1110 3222
rect -1322 3073 -1304 3189
rect -1124 3073 -1110 3189
rect 9272 3121 9286 3237
rect 9402 3196 9416 3237
rect 9402 3134 9534 3196
rect 9402 3121 9416 3134
rect 9272 3104 9416 3121
rect -1322 3036 -1110 3073
rect 11358 3084 11516 3134
rect 11358 3050 11381 3084
rect 11415 3050 11457 3084
rect 11491 3050 11516 3084
rect -4458 2952 -4344 3030
rect -4458 2856 -18 2952
rect 1742 2926 3604 2952
rect 5236 2926 6768 2952
rect 1702 2856 3614 2926
rect 5236 2856 6822 2926
rect 8472 2882 9828 2952
rect 8472 2856 9802 2882
rect -4458 2792 -4344 2856
rect 9300 2814 9586 2856
rect 9198 2644 9356 2672
rect 9198 2528 9218 2644
rect 9334 2528 9356 2644
rect 9198 2504 9356 2528
rect 9488 2272 9584 2298
rect 9622 2272 9764 2298
rect -4470 2134 -4356 2212
rect -4470 2038 -620 2134
rect -4470 1974 -4356 2038
rect -868 1272 -620 2038
rect 9488 1332 9764 2272
rect -868 1234 -708 1272
rect 570 1234 3302 1330
rect 7206 1303 10110 1332
rect 7206 1269 10020 1303
rect 10054 1269 10110 1303
rect 7206 1236 10110 1269
rect -4474 1008 -4360 1084
rect 3060 1082 3162 1104
rect 3060 1030 3086 1082
rect 3138 1030 3162 1082
rect -4474 912 -810 1008
rect 3060 1006 3162 1030
rect 8864 1082 9930 1112
rect 8864 1065 10014 1082
rect 8864 1031 8884 1065
rect 8918 1031 8956 1065
rect 8990 1031 10014 1065
rect 8864 1024 10014 1031
rect 8864 982 9006 1024
rect 11358 988 11516 3050
rect -4474 846 -4360 912
rect -1308 718 -1110 760
rect -1308 602 -1266 718
rect -1150 602 -1110 718
rect -906 738 -810 912
rect 840 918 960 948
rect 840 866 874 918
rect 926 866 960 918
rect 840 836 960 866
rect 9726 852 10016 912
rect 10688 904 11516 988
rect -906 642 -712 738
rect 570 642 3274 738
rect 7162 644 7758 740
rect -1308 590 -1110 602
rect -1308 562 -1112 590
rect -2002 482 -1688 522
rect -2002 480 -1969 482
rect -1725 480 -1688 482
rect -2002 374 -1974 480
rect -1724 374 -1688 480
rect -1208 454 -1112 562
rect 1558 538 1722 552
rect 1558 422 1587 538
rect 1703 422 1722 538
rect 1558 406 1722 422
rect -2002 366 -1969 374
rect -1725 366 -1688 374
rect -2002 330 -1688 366
rect -2010 50 -730 146
rect 570 50 3490 146
rect -4466 -110 -4352 -42
rect -2010 -110 -1914 50
rect -4466 -206 -1914 -110
rect -4466 -280 -4352 -206
rect 7590 -234 7758 644
rect 9726 186 9820 852
rect 9726 154 9912 186
rect 9726 38 9759 154
rect 9875 38 9912 154
rect 9726 10 9912 38
rect -1232 -512 7758 -234
rect -1222 -1050 -908 -512
rect 2808 -1026 3086 -512
rect 6804 -1006 7082 -512
<< via1 >>
rect -1304 3182 -1124 3189
rect -1304 3076 -1264 3182
rect -1264 3076 -1158 3182
rect -1158 3076 -1124 3182
rect -1304 3073 -1124 3076
rect 9286 3121 9402 3237
rect 9218 2640 9334 2644
rect 9218 2534 9224 2640
rect 9224 2534 9330 2640
rect 9330 2534 9334 2640
rect 9218 2528 9334 2534
rect 3086 1073 3138 1082
rect 3086 1039 3096 1073
rect 3096 1039 3130 1073
rect 3130 1039 3138 1073
rect 3086 1030 3138 1039
rect -1266 602 -1150 718
rect 874 910 926 918
rect 874 876 883 910
rect 883 876 917 910
rect 917 876 926 910
rect 874 866 926 876
rect -1969 480 -1725 482
rect -1969 374 -1725 480
rect 1587 534 1703 538
rect 1587 428 1594 534
rect 1594 428 1700 534
rect 1700 428 1703 534
rect 1587 422 1703 428
rect -1969 366 -1725 374
rect 9759 38 9875 154
<< metal2 >>
rect -1990 4022 -1694 4026
rect -4450 3972 -1694 4022
rect -4450 3836 -1953 3972
rect -1737 3836 -1694 3972
rect -4450 3786 -1694 3836
rect -4450 3784 -1696 3786
rect 8692 3254 9416 3256
rect 8692 3237 9418 3254
rect -1322 3197 -1108 3228
rect -1322 3189 -1280 3197
rect -1144 3189 -1108 3197
rect -1322 3073 -1304 3189
rect -1124 3073 -1108 3189
rect -1322 3061 -1280 3073
rect -1144 3061 -1108 3073
rect -1322 3034 -1108 3061
rect 8692 3121 9286 3237
rect 9402 3121 9418 3237
rect 8692 3102 9418 3121
rect 8692 3100 9416 3102
rect 8692 2672 8848 3100
rect -4460 2560 8848 2672
rect 9192 2656 9358 2674
rect 9192 2644 9247 2656
rect 9303 2644 9358 2656
rect -4460 2404 8850 2560
rect 9192 2528 9218 2644
rect 9334 2528 9358 2644
rect 9192 2520 9247 2528
rect 9303 2520 9358 2528
rect 9192 2502 9358 2520
rect -4470 1494 8716 1776
rect 3064 1082 3164 1494
rect 3064 1030 3086 1082
rect 3138 1030 3164 1082
rect 3064 1008 3164 1030
rect 830 918 1242 950
rect 830 866 874 918
rect 926 910 1242 918
rect 926 866 1244 910
rect 830 834 1244 866
rect -1310 728 -1108 764
rect -1310 592 -1280 728
rect -1144 592 -1108 728
rect -1310 558 -1108 592
rect -2012 528 -1824 530
rect -2012 495 -1678 528
rect -2012 482 -1957 495
rect -1741 482 -1678 495
rect -2012 366 -1969 482
rect -1725 366 -1678 482
rect -2012 359 -1957 366
rect -1741 359 -1678 366
rect -2012 326 -1678 359
rect 1046 396 1244 834
rect 1546 538 3266 596
rect 1546 422 1587 538
rect 1703 534 3266 538
rect 1703 484 3068 534
rect 8520 518 8716 1494
rect 10286 518 10386 714
rect 1703 422 1740 484
rect 1546 400 1740 422
rect 8520 418 10386 518
rect 8520 416 8716 418
rect -2012 324 -1824 326
rect 1046 312 1242 396
rect 1046 270 3060 312
rect 1046 198 3266 270
rect 9040 164 9214 166
rect 9040 104 9354 164
rect 9040 -32 9090 104
rect 9306 -32 9354 104
rect 9724 154 12028 188
rect 9724 38 9759 154
rect 9875 38 12028 154
rect 9724 10 12028 38
rect 9040 -86 9354 -32
rect 9040 -338 9350 -86
rect 9040 -544 10228 -338
rect -4128 -688 -3384 -596
rect -4128 -3170 -4036 -688
rect -3476 -1038 -3384 -688
rect -26 -704 806 -612
rect -3420 -3170 -3328 -2822
rect -4132 -3242 -3328 -3170
rect -4132 -3262 -3330 -3242
rect -24 -3276 68 -704
rect 714 -1014 806 -704
rect 4068 -700 4812 -608
rect 806 -3276 898 -2774
rect 4068 -3132 4160 -700
rect 4720 -1014 4812 -700
rect 4768 -3132 4860 -2774
rect 4066 -3200 4860 -3132
rect 4066 -3224 4858 -3200
rect -30 -3368 898 -3276
rect 9886 -3468 10228 -544
<< via2 >>
rect -1953 3836 -1737 3972
rect -1280 3189 -1144 3197
rect -1280 3073 -1144 3189
rect -1280 3061 -1144 3073
rect 9247 2644 9303 2656
rect 9247 2600 9303 2644
rect 9247 2528 9303 2576
rect 9247 2520 9303 2528
rect -1280 718 -1144 728
rect -1280 602 -1266 718
rect -1266 602 -1150 718
rect -1150 602 -1144 718
rect -1280 592 -1144 602
rect -1957 482 -1741 495
rect -1957 366 -1741 482
rect -1957 359 -1741 366
rect 9090 -32 9306 104
<< metal3 >>
rect -2004 3972 -1680 4060
rect -2004 3836 -1953 3972
rect -1737 3836 -1680 3972
rect -2004 495 -1680 3836
rect -1322 3197 -1108 3228
rect -1322 3061 -1280 3197
rect -1144 3061 -1108 3197
rect -1322 3034 -1108 3061
rect -1306 850 -1108 3034
rect -1308 820 -1108 850
rect 9096 2674 9256 2676
rect 9096 2672 9354 2674
rect 9096 2656 9358 2672
rect 9096 2600 9247 2656
rect 9303 2600 9358 2656
rect 9096 2576 9358 2600
rect 9096 2520 9247 2576
rect 9303 2520 9358 2576
rect -1308 728 -1110 820
rect -1308 592 -1280 728
rect -1144 592 -1110 728
rect -1308 562 -1110 592
rect -2004 359 -1957 495
rect -1741 359 -1680 495
rect -2004 332 -1680 359
rect 9096 158 9358 2520
rect 9042 156 9358 158
rect 9038 104 9366 156
rect 9038 -32 9090 104
rect 9306 -32 9366 104
rect 9038 -88 9366 -32
use Cap_295fF  Cap_295fF_0
timestamp 1607692587
transform 1 0 -3586 0 1 -2862
box -36 -56 3244 1928
use Cap_300fF  Cap_300fF_0
timestamp 1607692587
transform 1 0 500 0 1 -2850
box -200 -58 3244 1930
use ResTrial2  ResTrial2_2
timestamp 1607692587
transform 1 0 -148 0 1 -1922
box -78 -36 346 30
use Cap_305fF  Cap_305fF_0
timestamp 1607692587
transform 1 0 4622 0 1 -2850
box -200 -58 3244 1930
use ResTrial2  ResTrial2_1
timestamp 1607692587
transform 1 0 3950 0 1 -1910
box -78 -36 346 30
use ResTrial2  ResTrial2_0
timestamp 1607692587
transform 1 0 8094 0 1 -1910
box -78 -36 346 30
use PFD  PFD_0
timestamp 1607692587
transform 1 0 -868 0 1 50
box -340 0 1658 1280
use CP  CP_0
timestamp 1607692587
transform 1 0 3186 0 1 52
box 0 0 4134 1280
use MUX  MUX_0
timestamp 1607692587
transform 1 0 9956 0 1 612
box 0 -30 816 596
use /mnt/c/Users/LENOVO/Documents/PLL/Layout/new/FD  FD_2
timestamp 1607692587
transform -1 0 1782 0 1 2856
box 0 0 1880 640
use /mnt/c/Users/LENOVO/Documents/PLL/Layout/new/FD  FD_1
timestamp 1607692587
transform -1 0 5388 0 1 2856
box 0 0 1880 640
use /mnt/c/Users/LENOVO/Documents/PLL/Layout/new/FD  FD_0
timestamp 1607692587
transform -1 0 8552 0 1 2856
box 0 0 1880 640
use VCO  VCO_0
timestamp 1607692587
transform -1 0 11252 0 1 2220
box 0 0 1804 1280
<< labels >>
rlabel metal1 s -4450 3448 -4450 3448 4 VDD
port 1 nsew
rlabel metal1 s -4470 2092 -4470 2092 4 VDD
port 1 nsew
rlabel metal1 s -4458 2910 -4458 2910 4 GND
port 2 nsew
rlabel metal1 s -4474 964 -4474 964 4 GND
port 2 nsew
rlabel metal2 s -4460 2538 -4460 2538 4 ENb_VCO
port 3 nsew
rlabel metal2 s -4470 1634 -4470 1634 4 ENb_CP
port 4 nsew
rlabel metal2 s -4450 3902 -4450 3902 4 REF
port 5 nsew
rlabel metal2 s 10056 -3468 10056 -3468 4 CLK
port 6 nsew
rlabel metal2 s 12028 98 12028 98 4 VCO_IN
port 7 nsew
<< end >>
