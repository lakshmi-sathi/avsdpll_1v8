VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO /mnt/c/Users/LENOVO/Documents/PLL/Layout/VCO
  CLASS CORE ;
  FOREIGN /mnt/c/Users/LENOVO/Documents/PLL/Layout/VCO ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.020 BY 6.400 ;
  SITE unithddb1 ;
  PIN VCtrl
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.288000 ;
    PORT
      LAYER li1 ;
        RECT 0.070 4.190 0.800 4.390 ;
    END
  END VCtrl
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 0.150 9.020 0.320 ;
      LAYER mcon ;
        RECT 0.120 0.150 0.290 0.320 ;
        RECT 0.460 0.150 0.630 0.320 ;
        RECT 0.800 0.150 0.970 0.320 ;
        RECT 1.140 0.150 1.310 0.320 ;
        RECT 1.480 0.150 1.650 0.320 ;
        RECT 1.820 0.150 1.990 0.320 ;
        RECT 2.160 0.150 2.330 0.320 ;
        RECT 2.500 0.150 2.670 0.320 ;
        RECT 2.840 0.150 3.010 0.320 ;
        RECT 3.180 0.150 3.350 0.320 ;
        RECT 3.520 0.150 3.690 0.320 ;
        RECT 3.860 0.150 4.030 0.320 ;
        RECT 4.200 0.150 4.370 0.320 ;
        RECT 4.540 0.150 4.710 0.320 ;
        RECT 4.880 0.150 5.050 0.320 ;
        RECT 5.220 0.150 5.390 0.320 ;
        RECT 5.560 0.150 5.730 0.320 ;
        RECT 5.900 0.150 6.070 0.320 ;
        RECT 6.240 0.150 6.410 0.320 ;
        RECT 6.580 0.150 6.750 0.320 ;
        RECT 6.920 0.150 7.090 0.320 ;
        RECT 7.260 0.150 7.430 0.320 ;
        RECT 7.600 0.150 7.770 0.320 ;
        RECT 7.940 0.150 8.110 0.320 ;
        RECT 8.280 0.150 8.450 0.320 ;
        RECT 8.620 0.150 8.790 0.320 ;
      LAYER met1 ;
        RECT 0.000 0.000 9.020 0.480 ;
    END
    PORT
      LAYER nwell ;
        RECT 3.740 3.440 9.020 6.400 ;
        RECT 0.480 2.350 9.020 3.440 ;
      LAYER li1 ;
        RECT 0.000 6.050 9.020 6.220 ;
        RECT 6.460 5.270 6.800 6.050 ;
      LAYER mcon ;
        RECT 0.120 6.050 0.290 6.220 ;
        RECT 0.460 6.050 0.630 6.220 ;
        RECT 0.800 6.050 0.970 6.220 ;
        RECT 1.140 6.050 1.310 6.220 ;
        RECT 1.480 6.050 1.650 6.220 ;
        RECT 1.820 6.050 1.990 6.220 ;
        RECT 2.160 6.050 2.330 6.220 ;
        RECT 2.500 6.050 2.670 6.220 ;
        RECT 2.840 6.050 3.010 6.220 ;
        RECT 3.180 6.050 3.350 6.220 ;
        RECT 3.520 6.050 3.690 6.220 ;
        RECT 3.860 6.050 4.030 6.220 ;
        RECT 4.200 6.050 4.370 6.220 ;
        RECT 4.540 6.050 4.710 6.220 ;
        RECT 4.880 6.050 5.050 6.220 ;
        RECT 5.220 6.050 5.390 6.220 ;
        RECT 5.560 6.050 5.730 6.220 ;
        RECT 5.900 6.050 6.070 6.220 ;
        RECT 6.240 6.050 6.410 6.220 ;
        RECT 6.580 6.050 6.750 6.220 ;
        RECT 6.920 6.050 7.090 6.220 ;
        RECT 7.260 6.050 7.430 6.220 ;
        RECT 7.600 6.050 7.770 6.220 ;
        RECT 7.940 6.050 8.110 6.220 ;
        RECT 8.280 6.050 8.450 6.220 ;
        RECT 8.620 6.050 8.790 6.220 ;
      LAYER met1 ;
        RECT 0.000 5.920 9.020 6.400 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.690 5.230 0.860 5.460 ;
        RECT 0.690 5.060 2.090 5.230 ;
        RECT 0.690 4.780 3.370 5.060 ;
        RECT 0.690 4.620 0.860 4.780 ;
        RECT 1.390 4.740 3.370 4.780 ;
        RECT 1.390 4.460 2.090 4.740 ;
        RECT 2.710 4.490 3.370 4.740 ;
        RECT 1.190 4.290 2.270 4.460 ;
        RECT 2.710 3.990 3.380 4.490 ;
        RECT 2.720 3.700 3.370 3.990 ;
        RECT 8.170 1.330 8.340 1.870 ;
      LAYER mcon ;
        RECT 2.950 4.250 3.120 4.420 ;
        RECT 2.950 3.780 3.120 3.950 ;
        RECT 8.170 1.500 8.340 1.670 ;
      LAYER met1 ;
        RECT 2.720 4.490 3.370 4.500 ;
        RECT 2.710 3.450 3.380 4.490 ;
        RECT 0.050 2.970 9.020 3.450 ;
        RECT 8.710 1.730 8.910 2.970 ;
        RECT 8.110 1.440 8.910 1.730 ;
    END
  END GND
  PIN Clk_Out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.469800 ;
    PORT
      LAYER li1 ;
        RECT 8.610 2.310 8.780 3.610 ;
        RECT 8.610 2.080 9.020 2.310 ;
        RECT 8.610 1.330 8.780 2.080 ;
    END
  END Clk_Out
  PIN ENb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.063000 ;
    PORT
      LAYER li1 ;
        RECT 6.470 4.810 6.810 4.900 ;
        RECT 6.460 4.560 6.810 4.810 ;
      LAYER mcon ;
        RECT 6.550 4.630 6.720 4.800 ;
      LAYER met1 ;
        RECT 6.490 4.570 8.900 4.880 ;
    END
  END ENb
  OBS
      LAYER li1 ;
        RECT 0.250 4.620 0.420 5.460 ;
        RECT 4.300 5.250 5.220 5.360 ;
        RECT 5.470 5.250 5.640 5.450 ;
        RECT 4.300 5.040 5.640 5.250 ;
        RECT 4.720 4.840 5.640 5.040 ;
        RECT 5.470 4.610 5.640 4.840 ;
        RECT 5.910 4.540 6.110 5.490 ;
        RECT 7.100 5.270 8.580 5.690 ;
        RECT 8.170 5.130 8.580 5.270 ;
        RECT 5.850 4.410 6.110 4.540 ;
        RECT 3.930 4.240 6.110 4.410 ;
        RECT 7.150 4.090 7.320 4.760 ;
        RECT 0.210 3.770 2.280 4.020 ;
        RECT 3.930 3.800 5.010 3.970 ;
        RECT 0.210 1.270 0.580 3.770 ;
        RECT 4.150 3.440 4.740 3.800 ;
        RECT 6.430 3.740 7.320 4.090 ;
        RECT 5.830 3.440 7.320 3.740 ;
        RECT 1.150 3.120 7.320 3.440 ;
        RECT 1.150 2.530 1.320 3.120 ;
        RECT 1.590 2.280 1.760 2.950 ;
        RECT 2.150 2.530 2.320 3.120 ;
        RECT 2.590 2.280 2.760 2.950 ;
        RECT 3.150 2.530 3.320 3.120 ;
        RECT 3.590 2.280 3.760 2.950 ;
        RECT 4.150 2.530 4.320 3.120 ;
        RECT 4.590 2.280 4.760 2.950 ;
        RECT 5.150 2.530 5.320 3.120 ;
        RECT 5.590 2.280 5.760 2.950 ;
        RECT 6.150 2.530 6.320 3.120 ;
        RECT 6.590 2.280 6.760 2.950 ;
        RECT 7.150 2.530 7.320 3.120 ;
        RECT 7.590 2.340 7.760 4.760 ;
        RECT 8.170 4.400 8.470 5.130 ;
        RECT 8.170 2.530 8.340 4.400 ;
        RECT 0.820 2.110 1.420 2.280 ;
        RECT 1.590 2.110 2.420 2.280 ;
        RECT 2.590 2.110 3.420 2.280 ;
        RECT 3.590 2.110 4.420 2.280 ;
        RECT 4.590 2.110 5.420 2.280 ;
        RECT 5.590 2.110 6.420 2.280 ;
        RECT 6.590 2.110 7.420 2.280 ;
        RECT 1.150 1.270 1.320 1.860 ;
        RECT 1.590 1.440 1.760 2.110 ;
        RECT 2.150 1.270 2.320 1.860 ;
        RECT 2.590 1.440 2.760 2.110 ;
        RECT 3.150 1.270 3.320 1.860 ;
        RECT 3.590 1.440 3.760 2.110 ;
        RECT 4.150 1.270 4.320 1.860 ;
        RECT 4.590 1.440 4.760 2.110 ;
        RECT 5.150 1.270 5.320 1.860 ;
        RECT 5.590 1.440 5.760 2.110 ;
        RECT 6.150 1.270 6.320 1.860 ;
        RECT 6.590 1.440 6.760 2.110 ;
        RECT 7.590 2.050 8.430 2.340 ;
        RECT 7.150 1.330 7.320 1.860 ;
        RECT 7.000 1.270 7.320 1.330 ;
        RECT 0.210 0.950 7.320 1.270 ;
        RECT 7.000 0.900 7.320 0.950 ;
        RECT 7.150 0.770 7.320 0.900 ;
        RECT 7.590 0.770 7.760 2.050 ;
      LAYER mcon ;
        RECT 0.250 5.060 0.420 5.230 ;
        RECT 4.360 5.100 4.580 5.300 ;
        RECT 5.910 5.120 6.080 5.290 ;
        RECT 7.110 5.390 7.280 5.560 ;
        RECT 7.920 2.110 8.090 2.280 ;
      LAYER met1 ;
        RECT 4.330 5.310 4.640 5.360 ;
        RECT 7.050 5.340 7.340 5.620 ;
        RECT 0.190 5.000 4.640 5.310 ;
        RECT 5.850 5.070 7.350 5.340 ;
        RECT 0.760 2.060 8.130 2.340 ;
        RECT 0.760 2.050 8.120 2.060 ;
  END
END /mnt/c/Users/LENOVO/Documents/PLL/Layout/VCO
END LIBRARY

