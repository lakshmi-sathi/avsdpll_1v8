magic
tech sky130A
timestamp 1605269755
<< nwell >>
rect -59 287 416 392
rect -11 231 416 287
rect 235 180 416 231
rect 249 128 416 180
rect 249 -90 551 128
rect 249 -91 508 -90
rect 249 -167 366 -91
<< nmos >>
rect 455 265 503 280
rect 455 214 491 229
rect 0 146 84 161
rect 0 90 180 105
rect 0 33 36 48
rect 51 -156 66 -120
rect 108 -156 123 24
rect 164 -156 179 -72
rect 431 -165 446 -129
rect 482 -177 497 -129
<< pmos >>
rect 7 282 72 297
rect 139 282 204 297
rect 285 265 381 280
rect 285 214 357 229
rect 300 -17 315 48
rect 431 -31 446 41
rect 482 -55 497 41
rect 300 -149 315 -84
<< ndiff >>
rect 455 305 503 309
rect 455 288 470 305
rect 487 288 503 305
rect 455 280 503 288
rect 0 186 84 194
rect 0 169 29 186
rect 46 169 63 186
rect 80 169 84 186
rect 0 161 84 169
rect 455 259 503 265
rect 455 242 479 259
rect 496 242 503 259
rect 455 238 503 242
rect 455 229 491 238
rect 455 206 491 214
rect 455 189 465 206
rect 482 189 491 206
rect 455 183 491 189
rect 0 138 84 146
rect 0 130 180 138
rect 0 113 4 130
rect 21 113 38 130
rect 55 113 72 130
rect 89 113 106 130
rect 123 113 140 130
rect 157 113 180 130
rect 0 105 180 113
rect 0 57 180 90
rect 0 48 36 57
rect 0 25 36 33
rect 0 8 10 25
rect 27 8 36 25
rect 0 0 36 8
rect 75 -120 108 24
rect 18 -130 51 -120
rect 18 -147 26 -130
rect 43 -147 51 -130
rect 18 -156 51 -147
rect 66 -156 108 -120
rect 123 1 156 24
rect 123 -16 131 1
rect 148 -16 156 1
rect 123 -33 156 -16
rect 123 -50 131 -33
rect 148 -50 156 -33
rect 123 -67 156 -50
rect 123 -84 131 -67
rect 148 -72 156 -67
rect 148 -84 164 -72
rect 123 -101 164 -84
rect 123 -118 131 -101
rect 148 -118 164 -101
rect 123 -135 164 -118
rect 123 -152 131 -135
rect 148 -152 164 -135
rect 123 -156 164 -152
rect 179 -76 212 -72
rect 179 -93 187 -76
rect 204 -93 212 -76
rect 179 -110 212 -93
rect 179 -127 187 -110
rect 204 -127 212 -110
rect 179 -156 212 -127
rect 400 -139 431 -129
rect 400 -156 406 -139
rect 423 -156 431 -139
rect 400 -165 431 -156
rect 446 -153 482 -129
rect 446 -165 459 -153
rect 455 -170 459 -165
rect 476 -170 482 -153
rect 455 -177 482 -170
rect 497 -144 526 -129
rect 497 -161 505 -144
rect 522 -161 526 -144
rect 497 -177 526 -161
<< pdiff >>
rect 7 322 72 330
rect 7 305 11 322
rect 28 305 45 322
rect 62 305 72 322
rect 139 322 204 330
rect 7 297 72 305
rect 7 274 72 282
rect 7 257 15 274
rect 32 257 51 274
rect 68 257 72 274
rect 139 305 143 322
rect 160 305 177 322
rect 194 305 204 322
rect 139 297 204 305
rect 285 304 381 310
rect 285 287 289 304
rect 306 287 323 304
rect 340 287 381 304
rect 139 274 204 282
rect 285 280 381 287
rect 7 249 72 257
rect 139 257 148 274
rect 165 257 182 274
rect 199 257 204 274
rect 139 249 204 257
rect 285 259 381 265
rect 285 242 289 259
rect 306 242 323 259
rect 340 242 381 259
rect 285 238 381 242
rect 285 229 357 238
rect 285 206 357 214
rect 285 189 289 206
rect 306 189 323 206
rect 340 189 357 206
rect 285 183 357 189
rect 267 43 300 48
rect 267 26 275 43
rect 292 26 300 43
rect 267 9 300 26
rect 267 -8 275 9
rect 292 -8 300 9
rect 267 -17 300 -8
rect 315 38 348 48
rect 315 21 323 38
rect 340 21 348 38
rect 315 4 348 21
rect 315 -13 323 4
rect 340 -13 348 4
rect 315 -17 348 -13
rect 400 37 431 41
rect 400 20 406 37
rect 423 20 431 37
rect 400 3 431 20
rect 400 -14 406 3
rect 423 -14 431 3
rect 400 -31 431 -14
rect 446 37 482 41
rect 446 20 459 37
rect 476 20 482 37
rect 446 3 482 20
rect 446 -14 459 3
rect 476 -14 482 3
rect 446 -31 482 -14
rect 455 -55 482 -31
rect 497 37 527 41
rect 497 20 504 37
rect 521 20 527 37
rect 497 3 527 20
rect 497 -14 504 3
rect 521 -14 527 3
rect 497 -55 527 -14
rect 267 -88 300 -84
rect 267 -105 275 -88
rect 292 -105 300 -88
rect 267 -124 300 -105
rect 267 -141 275 -124
rect 292 -141 300 -124
rect 267 -149 300 -141
rect 315 -94 348 -84
rect 315 -111 323 -94
rect 340 -111 348 -94
rect 315 -128 348 -111
rect 315 -145 323 -128
rect 340 -145 348 -128
rect 315 -149 348 -145
<< ndiffc >>
rect 470 288 487 305
rect 29 169 46 186
rect 63 169 80 186
rect 479 242 496 259
rect 465 189 482 206
rect 4 113 21 130
rect 38 113 55 130
rect 72 113 89 130
rect 106 113 123 130
rect 140 113 157 130
rect 10 8 27 25
rect 26 -147 43 -130
rect 131 -16 148 1
rect 131 -50 148 -33
rect 131 -84 148 -67
rect 131 -118 148 -101
rect 131 -152 148 -135
rect 187 -93 204 -76
rect 187 -127 204 -110
rect 406 -156 423 -139
rect 459 -170 476 -153
rect 505 -161 522 -144
<< pdiffc >>
rect 11 305 28 322
rect 45 305 62 322
rect 15 257 32 274
rect 51 257 68 274
rect 143 305 160 322
rect 177 305 194 322
rect 289 287 306 304
rect 323 287 340 304
rect 148 257 165 274
rect 182 257 199 274
rect 289 242 306 259
rect 323 242 340 259
rect 289 189 306 206
rect 323 189 340 206
rect 275 26 292 43
rect 275 -8 292 9
rect 323 21 340 38
rect 323 -13 340 4
rect 406 20 423 37
rect 406 -14 423 3
rect 459 20 476 37
rect 459 -14 476 3
rect 504 20 521 37
rect 504 -14 521 3
rect 275 -105 292 -88
rect 275 -141 292 -124
rect 323 -111 340 -94
rect 323 -145 340 -128
<< psubdiff >>
rect 531 289 548 301
rect 531 260 548 272
rect 531 221 548 233
rect 531 192 548 204
rect -2 -44 10 -27
rect 27 -44 39 -27
rect -67 -233 -55 -216
rect -38 -233 -25 -216
rect 17 -233 29 -216
rect 46 -233 59 -216
rect 101 -233 113 -216
rect 130 -233 143 -216
rect 185 -234 197 -217
rect 214 -234 227 -217
rect 269 -234 281 -217
rect 298 -234 311 -217
rect 409 -222 421 -205
rect 438 -222 450 -205
rect 477 -222 489 -205
rect 506 -222 518 -205
<< nsubdiff >>
rect -32 357 -20 374
rect -3 357 9 374
rect 50 357 62 374
rect 79 357 91 374
rect 132 357 144 374
rect 161 357 173 374
rect 214 357 226 374
rect 243 357 255 374
rect 296 357 308 374
rect 325 357 337 374
rect 302 113 346 117
rect 302 93 314 113
rect 334 93 346 113
rect 302 89 346 93
<< psubdiffcont >>
rect 531 272 548 289
rect 531 204 548 221
rect 10 -44 27 -27
rect -55 -233 -38 -216
rect 29 -233 46 -216
rect 113 -233 130 -216
rect 197 -234 214 -217
rect 281 -234 298 -217
rect 421 -222 438 -205
rect 489 -222 506 -205
<< nsubdiffcont >>
rect -20 357 -3 374
rect 62 357 79 374
rect 144 357 161 374
rect 226 357 243 374
rect 308 357 325 374
rect 314 93 334 113
<< poly >>
rect 92 298 119 306
rect 92 297 97 298
rect -6 282 7 297
rect 72 282 97 297
rect 92 281 97 282
rect 114 297 119 298
rect 114 282 139 297
rect 204 282 217 297
rect 114 281 119 282
rect 92 273 119 281
rect 97 161 114 273
rect 272 265 285 280
rect 381 273 455 280
rect 381 265 407 273
rect 391 262 407 265
rect 398 256 407 262
rect 424 265 455 273
rect 503 265 516 280
rect 424 262 438 265
rect 424 256 432 262
rect 398 251 432 256
rect 272 214 285 229
rect 357 223 455 229
rect 357 214 402 223
rect 397 206 402 214
rect 419 214 455 223
rect 491 214 506 229
rect 419 206 424 214
rect 397 201 424 206
rect 402 198 419 201
rect -24 146 0 161
rect 84 146 114 161
rect -24 105 -9 146
rect -62 92 0 105
rect -62 75 -57 92
rect -40 90 0 92
rect 180 90 193 105
rect -40 75 -35 90
rect -62 67 -35 75
rect 55 48 207 49
rect 300 48 315 61
rect -13 33 0 48
rect 36 38 207 48
rect 36 33 182 38
rect 108 24 123 33
rect 28 -80 66 -75
rect 28 -97 36 -80
rect 53 -97 66 -80
rect 28 -102 66 -97
rect 51 -120 66 -102
rect 171 21 182 33
rect 199 21 207 38
rect 171 16 207 21
rect 431 41 446 54
rect 482 41 497 54
rect 300 -37 315 -17
rect 291 -42 324 -37
rect 164 -59 299 -42
rect 316 -59 324 -42
rect 164 -72 179 -59
rect 291 -64 324 -59
rect 300 -84 315 -64
rect 431 -71 446 -31
rect 482 -65 497 -55
rect 418 -76 446 -71
rect 479 -72 497 -65
rect 415 -93 423 -76
rect 440 -93 447 -76
rect 468 -81 497 -72
rect 418 -98 446 -93
rect 431 -129 446 -98
rect 468 -98 473 -81
rect 490 -98 497 -81
rect 468 -106 497 -98
rect 479 -112 497 -106
rect 482 -129 497 -112
rect 51 -171 66 -156
rect 108 -165 123 -156
rect 164 -165 179 -156
rect 300 -162 315 -149
rect 108 -180 179 -165
rect 431 -180 446 -165
rect 482 -190 497 -177
<< polycont >>
rect 97 281 114 298
rect 407 256 424 273
rect 402 206 419 223
rect -57 75 -40 92
rect 36 -97 53 -80
rect 182 21 199 38
rect 299 -59 316 -42
rect 423 -93 440 -76
rect 473 -98 490 -81
<< locali >>
rect -85 374 555 392
rect -85 357 -20 374
rect -3 357 62 374
rect 79 357 144 374
rect 161 357 226 374
rect 243 357 308 374
rect 325 357 555 374
rect -85 344 555 357
rect 17 324 59 344
rect 3 322 74 324
rect 3 305 11 322
rect 28 305 45 322
rect 62 305 74 322
rect 3 303 74 305
rect 94 322 204 323
rect 94 305 143 322
rect 160 305 177 322
rect 194 305 204 322
rect 94 304 204 305
rect 94 298 117 304
rect 94 281 97 298
rect 114 281 117 298
rect 237 293 262 344
rect 285 305 503 316
rect 7 274 76 276
rect 7 257 15 274
rect 32 257 51 274
rect 68 257 76 274
rect 94 273 117 281
rect 139 274 207 275
rect 7 256 76 257
rect 139 257 148 274
rect 165 257 182 274
rect 199 257 207 274
rect 139 256 207 257
rect 236 260 262 293
rect 281 304 470 305
rect 281 287 289 304
rect 306 287 323 304
rect 340 299 470 304
rect 340 287 381 299
rect 455 288 470 299
rect 487 288 503 305
rect 455 286 503 288
rect 526 289 554 306
rect 398 270 407 273
rect 236 259 351 260
rect -33 230 76 256
rect -33 144 -6 230
rect 150 194 194 256
rect 236 242 289 259
rect 306 242 323 259
rect 340 242 351 259
rect 236 237 351 242
rect 368 256 407 270
rect 424 268 432 273
rect 526 272 531 289
rect 548 272 554 289
rect 424 256 453 268
rect 526 263 554 272
rect 519 260 554 263
rect 368 251 453 256
rect 368 208 385 251
rect 427 250 453 251
rect 281 206 385 208
rect 211 194 248 195
rect 17 186 248 194
rect 281 189 289 206
rect 306 189 323 206
rect 340 189 385 206
rect 281 186 385 189
rect 402 223 419 231
rect 17 169 29 186
rect 46 169 63 186
rect 80 169 248 186
rect 402 169 419 206
rect 436 207 453 250
rect 471 259 554 260
rect 471 242 479 259
rect 496 242 554 259
rect 471 238 554 242
rect 519 234 554 238
rect 526 221 554 234
rect 436 206 491 207
rect 436 189 465 206
rect 482 189 491 206
rect 436 185 491 189
rect 526 204 531 221
rect 548 204 554 221
rect 526 184 554 204
rect 17 168 419 169
rect -33 137 7 144
rect 211 139 419 168
rect -33 131 27 137
rect -33 130 180 131
rect -33 118 4 130
rect -22 113 4 118
rect 21 113 38 130
rect 55 113 72 130
rect 89 113 106 130
rect 123 113 140 130
rect 157 113 180 130
rect -22 112 180 113
rect 302 113 481 117
rect -66 92 -39 100
rect -66 75 -57 92
rect -40 75 -39 92
rect 302 93 314 113
rect 334 93 481 113
rect 302 87 481 93
rect -66 -76 -39 75
rect 454 83 481 87
rect 174 38 207 48
rect 274 43 293 51
rect 274 38 275 43
rect 8 25 29 27
rect 0 8 10 25
rect 27 8 36 25
rect 8 -24 29 8
rect 130 1 149 24
rect 174 21 182 38
rect 199 21 207 38
rect 225 26 275 38
rect 292 26 293 43
rect 225 9 293 26
rect 225 3 275 9
rect 130 -16 131 1
rect 148 -16 149 1
rect 1 -27 37 -24
rect 1 -44 10 -27
rect 27 -44 37 -27
rect 1 -47 37 -44
rect 130 -33 149 -16
rect 130 -50 131 -33
rect 148 -50 149 -33
rect 130 -67 149 -50
rect -15 -76 62 -74
rect -66 -80 62 -76
rect -66 -97 36 -80
rect 53 -97 62 -80
rect -66 -103 62 -97
rect 130 -84 131 -67
rect 148 -84 149 -67
rect 187 -6 275 3
rect 187 -8 246 -6
rect 187 -25 195 -8
rect 212 -22 246 -8
rect 274 -8 275 -6
rect 292 -8 293 9
rect 274 -17 293 -8
rect 322 38 341 48
rect 322 21 323 38
rect 340 21 341 38
rect 322 4 341 21
rect 322 -13 323 4
rect 340 -13 341 4
rect 212 -25 216 -22
rect 187 -28 216 -25
rect 187 -72 212 -28
rect 322 -39 341 -13
rect 291 -42 341 -39
rect 291 -59 299 -42
rect 316 -59 341 -42
rect 403 37 425 45
rect 403 20 406 37
rect 423 20 425 37
rect 403 3 425 20
rect 403 -14 406 3
rect 423 -14 425 3
rect 403 -42 425 -14
rect 454 37 477 83
rect 454 20 459 37
rect 476 20 477 37
rect 454 3 477 20
rect 454 -14 459 3
rect 476 -14 477 3
rect 454 -25 477 -14
rect 504 41 522 45
rect 504 37 533 41
rect 521 20 533 37
rect 504 3 533 20
rect 521 -14 533 3
rect 403 -59 487 -42
rect 504 -55 533 -14
rect 291 -62 341 -59
rect 130 -101 149 -84
rect -66 -105 2 -103
rect 25 -130 43 -120
rect 25 -147 26 -130
rect 25 -170 43 -147
rect 130 -124 131 -101
rect 148 -124 149 -101
rect 130 -135 149 -124
rect 130 -152 131 -135
rect 148 -152 149 -135
rect 186 -76 212 -72
rect 468 -72 487 -59
rect 186 -93 187 -76
rect 204 -93 212 -76
rect 186 -110 212 -93
rect 186 -127 187 -110
rect 204 -127 212 -110
rect 186 -139 212 -127
rect 248 -88 294 -80
rect 248 -105 275 -88
rect 292 -105 294 -88
rect 248 -107 294 -105
rect 248 -124 261 -107
rect 278 -124 294 -107
rect 248 -141 275 -124
rect 292 -141 294 -124
rect 248 -149 294 -141
rect 321 -94 342 -82
rect 366 -93 372 -76
rect 389 -93 423 -76
rect 440 -93 448 -76
rect 468 -81 490 -72
rect 321 -124 323 -94
rect 340 -124 342 -94
rect 468 -98 473 -81
rect 468 -101 490 -98
rect 467 -106 490 -101
rect 467 -110 485 -106
rect 321 -128 342 -124
rect 321 -145 323 -128
rect 340 -145 342 -128
rect 130 -162 149 -152
rect 321 -153 342 -145
rect 402 -127 485 -110
rect 402 -139 424 -127
rect 516 -129 533 -55
rect 402 -156 406 -139
rect 423 -156 424 -139
rect 503 -144 533 -129
rect 402 -165 424 -156
rect 455 -153 477 -145
rect 15 -192 43 -170
rect 8 -200 43 -192
rect 455 -170 459 -153
rect 476 -170 477 -153
rect 455 -193 477 -170
rect 503 -161 505 -144
rect 522 -161 533 -144
rect 503 -177 533 -161
rect 451 -200 480 -193
rect -85 -205 555 -200
rect -85 -216 421 -205
rect -85 -233 -55 -216
rect -38 -233 29 -216
rect 46 -233 113 -216
rect 130 -217 421 -216
rect 130 -233 197 -217
rect -85 -234 197 -233
rect 214 -234 281 -217
rect 298 -222 421 -217
rect 438 -222 489 -205
rect 506 -222 555 -205
rect 298 -234 555 -222
rect -85 -248 555 -234
<< viali >>
rect 314 93 334 113
rect 195 -25 212 -8
rect 131 -118 148 -107
rect 131 -124 148 -118
rect 261 -124 278 -107
rect 372 -93 389 -76
rect 323 -111 340 -107
rect 323 -124 340 -111
<< metal1 >>
rect 303 113 348 126
rect 303 93 314 113
rect 334 93 348 113
rect 303 81 348 93
rect 186 -2 221 1
rect 186 -31 189 -2
rect 218 -31 221 -2
rect 317 -5 348 81
rect 186 -34 221 -31
rect 30 -103 59 -74
rect 125 -107 284 -101
rect 125 -124 131 -107
rect 148 -124 261 -107
rect 278 -124 284 -107
rect 125 -130 284 -124
rect 317 -107 348 -31
rect 365 -72 397 -69
rect 365 -98 368 -72
rect 394 -98 397 -72
rect 365 -101 397 -98
rect 317 -124 323 -107
rect 340 -124 348 -107
rect 317 -130 348 -124
<< via1 >>
rect 189 -8 218 -2
rect 189 -25 195 -8
rect 195 -25 212 -8
rect 212 -25 218 -8
rect 189 -31 218 -25
rect 368 -76 394 -72
rect 368 -93 372 -76
rect 372 -93 389 -76
rect 389 -93 394 -76
rect 368 -98 394 -93
<< metal2 >>
rect 186 -2 221 1
rect 186 -31 189 -2
rect 218 -29 392 -2
rect 218 -31 221 -29
rect 186 -34 221 -31
rect 366 -69 392 -29
rect 365 -72 397 -69
rect 365 -98 368 -72
rect 394 -98 397 -72
rect 365 -101 397 -98
<< labels >>
rlabel locali -61 -104 -34 -77 1 Clk_Ref
port 3 n
rlabel locali 182 26 199 43 1 Clk2
port 4 n
rlabel locali -85 344 -85 392 3 VDD
port 5 e
rlabel locali -85 -248 -85 -200 3 GND
port 6 e
rlabel locali 409 299 426 316 1 Up
port 7 n
rlabel locali 516 -99 533 -82 1 Down
port 8 n
<< end >>
