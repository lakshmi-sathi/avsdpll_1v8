*---------PLL---------
.include sky130nm.lib

xx1 clk_ref clk_vco_by_8 up down phase_detector
xx2 up down vin_vco chpmp
xx3 vin_vco clk_out vcoscillator

xx5 clk_out 4 freqdiv2
xx6 4 3 freqdiv2
x7 3 clk_vco_by_8 freqdiv2
c3 clk_vco_by_8 0 1f

v1 clk_ref 0 PULSE 0 1.8 10p 60p 60p 100ns 200ns
v2 1 0 1.8

*PD-----------------
.subckt phase_detector clk1 clk2 up down
xm1 1 clk1 3 1 sky130_fd_pr__pfet_01v8 l=150n w=420n 
xm2 3 clk1 4 0 sky130_fd_pr__nfet_01v8 l=150n w=420n
xm3 4 clk2 0 0 sky130_fd_pr__nfet_01v8 l=150n w=420n

xm4 1 clk2 6 1 sky130_fd_pr__pfet_01v8 l=150n w=420n 
xm5 6 clk2 7 0 sky130_fd_pr__nfet_01v8 l=150n w=420n
xm6 7 clk1 0 0 sky130_fd_pr__nfet_01v8 l=150n w=420n

xm7 8 clk1 3 0 sky130_fd_pr__nfet_01v8 l=150n w=1440n 
xm8 clk1 clk1 8 1 sky130_fd_pr__pfet_01v8 l=150n w=1440n

xm9 9 clk2 6 0 sky130_fd_pr__nfet_01v8 l=150n w=1440n
xm10 clk2 clk2 9 1 sky130_fd_pr__pfet_01v8 l=150n w=1440n

*output cap
c1 8 0 0.9f
c2 9 0 0.9f

*buffer
xm11 1 8 10 1 sky130_fd_pr__pfet_01v8 l=150n w=720n 
xm12 10 8 0 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm15 1 10 up 1 sky130_fd_pr__pfet_01v8 l=150n w=1080n 
xm16 up 10 0 0 sky130_fd_pr__nfet_01v8 l=150n w=540n
xm13 1 9 11 1 sky130_fd_pr__pfet_01v8 l=150n w=720n 
xm17 11 9 0 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm18 1 11 down 1 sky130_fd_pr__pfet_01v8 l=150n w=1080n
xm14 down 11 0 0 sky130_fd_pr__nfet_01v8 l=150n w=540n

v1 1 0 1.8

.ends phase_detector
*--------------------

*ChargePump---------------
.subckt chpmp up down out
*---Top 2---
xm1 2 0 1 1 sky130_fd_pr__pfet_01v8 l=150n w=840n 
xm2 4 up 1 1 sky130_fd_pr__pfet_01v8 l=150n w=420n
*---Left Top SC Transistor--- 
xm3 5 3 2 1 sky130_fd_pr__pfet_01v8 l=600n w=2400n 
xm4 3 3 5 7 sky130_fd_pr__pfet_01v8 l=150n w=9600n  
*---Right Top SC Transistor---
xm5 6 3 4 1 sky130_fd_pr__pfet_01v8 l=600n w=1200n 
xm6 out 3 6 7 sky130_fd_pr__pfet_01v8 l=150n w=4800n


*---Right Bottom SC Transistor---
xm7 out 8 10 15 sky130_fd_pr__nfet_01v8 l=150n w=4800n
xm8 10 8 11 0 sky130_fd_pr__nfet_01v8 l=600n w=1200n
*---Left Bottom SC Transistor---
xm9 9 8 3 15 sky130_fd_pr__nfet_01v8 l=150n w=9600n
xm10 12 8 9 0 sky130_fd_pr__nfet_01v8 l=600n w=2400n
*---Bottom 2---
xm11 0 1 12 0 sky130_fd_pr__nfet_01v8 l=150n w=420n
xm12 0 down 11 0 sky130_fd_pr__nfet_01v8 l=150n w=420n

*---Current Source---
xm16 16 16 0 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm17 8 16 16 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
*---Mirroring Iref-----
xm13 13 8 8 15 sky130_fd_pr__nfet_01v8 l=150n w=2400n
xm14 14 8 13 0 sky130_fd_pr__nfet_01v8 l=600n w=600n
xm15 0 1 14 0 sky130_fd_pr__nfet_01v8 l=150n w=420n


r1 15 16 480

c1 out 0 0.52f
v1 1 0 1.8
v2 7 0 1.4 
v3 15 0 0.4
.ends chpmp
*------------------

*LPF----------------
c1 vin_vco 0 0.2f
c2 5 0 1f
r1 vin_vco 5 10
*-------------------

*VCO----------------
.subckt vcoscillator vin vout
xm1 vp vn 0 0 sky130_fd_pr__nfet_01v8 l=200n w=400n
xm2 vp vp 1 1 sky130_fd_pr__pfet_01v8 l=200n w=2000n
r1 vn vin 1
*xu1 osc_fb Osc inv_20_10
xm3 1 osc_fb vout 1 sky130_fd_pr__pfet_01v8 l=150n w=2400n 
xm4 vout osc_fb 0 0 sky130_fd_pr__nfet_01v8 l=150n w=1200n
xx1 7 osc_fb vp vn cs_inv
xx2 6 7 vp vn cs_inv
xx3 5 6 vp vn cs_inv
xx4 4 5 vp vn cs_inv
xx5 3 4 vp vn cs_inv
xx6 2 3 vp vn cs_inv
xx7 osc_fb 2 vp vn cs_inv
c1 vout 0 0.1f

v1 1 0 1.8
.ends vcoscillator

.subckt cs_inv in out vp vn
xm1 3 vn 0 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm2 2 vp 1 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm3 out in 2 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm4 out in 3 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

c1 out 0 1f
v1 1 0 1.8
.ends cs_inv
*----------------------

**VCO---------------------
*.subckt vcoscillator vin vout
*xm1 10 vout 3 10 sky130_fd_pr__pfet_01v8 l=150n w=900n
*xm2 3 vout 9 9  sky130_fd_pr__nfet_01v8 l=150n w=360n
*
*xm3 10 3 4 10 sky130_fd_pr__pfet_01v8 l=150n w=900n
*xm4 4 3 9 9 sky130_fd_pr__nfet_01v8 l=150n w=360n
*
*xm5 10 4 vout 10 sky130_fd_pr__pfet_01v8 l=150n w=900n
*xm6 vout 4 9 9 sky130_fd_pr__nfet_01v8 l=150n w=360n
*
*xm7 10 5 1 1 sky130_fd_pr__pfet_01v8 l=150n w=420n
*xm8 5 5 1 1 sky130_fd_pr__pfet_01v8 l=150n w=420n
*xm9 5 vin 0 0 sky130_fd_pr__nfet_01v8 l=150n w=2400n
*xm10 9 vin 0 0 sky130_fd_pr__nfet_01v8 l=150n w=2400n
*
*c1 2 0 0.1f
*v1 1 0 1.8
*.ends vcoscillator
**--------------------------

*FreqDiv by 2-----------
.subckt freqdiv2 clkin clkout 
xm1 1 5 2 1 sky130_fd_pr__pfet_01v8 l=150n w=3050n 
xm2 2 clkin 0 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm3 1 2 4 1 sky130_fd_pr__pfet_01v8 l=150n w=420n 
xm4 4 clkin 0 0 sky130_fd_pr__nfet_01v8 l=150n w=840n

xm5 1 clkin 5 1 sky130_fd_pr__pfet_01v8 l=150n w=420n 
xm6 5 4 0 0 sky130_fd_pr__nfet_01v8 l=150n w=840n

c1 5 0 0.8f

xm7 1 5 6 1 sky130_fd_pr__pfet_01v8 l=150n w=900n 
xm8 6 5 0 0 sky130_fd_pr__nfet_01v8 l=150n w=450n

xm9 1 6 clkout 1 sky130_fd_pr__pfet_01v8 l=150n w=900n 
xm10 clkout 6 0 0 sky130_fd_pr__nfet_01v8 l=150n w=450n


v1 1 0 1.8
.ends freqdiv2
*-----------------------


*simulation
.ic V(vin_vco) = 0
.control
tran 1ns 40us
plot v(up)+8 v(down)+6 v(clk_ref)+4 v(vin_vco)+2  v(clk_out) 
.endc
.end 
