VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO CP
  CLASS CORE ;
  FOREIGN CP ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.670 BY 6.400 ;
  SITE unithddb1 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.120 4.670 20.660 6.260 ;
        RECT 0.120 4.360 8.160 4.670 ;
        RECT 1.960 4.230 8.160 4.360 ;
        RECT 2.300 4.080 8.160 4.230 ;
        RECT 2.410 4.030 8.160 4.080 ;
        RECT 11.580 3.930 20.660 4.670 ;
        RECT 11.580 3.890 19.420 3.930 ;
        RECT 11.580 3.880 12.880 3.890 ;
        RECT 11.580 3.580 12.510 3.880 ;
      LAYER li1 ;
        RECT 0.000 6.070 20.660 6.240 ;
        RECT 2.480 5.850 20.480 6.070 ;
        RECT 13.380 4.200 20.150 4.410 ;
      LAYER mcon ;
        RECT 0.210 6.070 0.380 6.240 ;
        RECT 0.550 6.070 0.720 6.240 ;
        RECT 0.890 6.070 1.060 6.240 ;
        RECT 1.230 6.070 1.400 6.240 ;
        RECT 1.570 6.070 1.740 6.240 ;
        RECT 1.910 6.070 2.080 6.240 ;
        RECT 2.250 6.070 2.420 6.240 ;
        RECT 2.590 6.070 2.760 6.240 ;
        RECT 2.930 6.070 3.100 6.240 ;
        RECT 3.270 6.070 3.440 6.240 ;
        RECT 3.610 6.070 3.780 6.240 ;
        RECT 3.950 6.070 4.120 6.240 ;
        RECT 4.290 6.070 4.460 6.240 ;
        RECT 4.630 6.070 4.800 6.240 ;
        RECT 4.970 6.070 5.140 6.240 ;
        RECT 5.310 6.070 5.480 6.240 ;
        RECT 5.650 6.070 5.820 6.240 ;
        RECT 5.990 6.070 6.160 6.240 ;
        RECT 6.330 6.070 6.500 6.240 ;
        RECT 6.670 6.070 6.840 6.240 ;
        RECT 7.010 6.070 7.180 6.240 ;
        RECT 7.350 6.070 7.520 6.240 ;
        RECT 7.690 6.070 7.860 6.240 ;
        RECT 8.030 6.070 8.200 6.240 ;
        RECT 8.370 6.070 8.540 6.240 ;
        RECT 8.710 6.070 8.880 6.240 ;
        RECT 9.050 6.070 9.220 6.240 ;
        RECT 9.390 6.070 9.560 6.240 ;
        RECT 9.730 6.070 9.900 6.240 ;
        RECT 10.070 6.070 10.240 6.240 ;
        RECT 10.410 6.070 10.580 6.240 ;
        RECT 10.750 6.070 10.920 6.240 ;
        RECT 11.090 6.070 11.260 6.240 ;
        RECT 11.430 6.070 11.600 6.240 ;
        RECT 11.770 6.070 11.940 6.240 ;
        RECT 12.110 6.070 12.280 6.240 ;
        RECT 12.450 6.070 12.620 6.240 ;
        RECT 12.790 6.070 12.960 6.240 ;
        RECT 13.130 6.070 13.300 6.240 ;
        RECT 13.470 6.070 13.640 6.240 ;
        RECT 13.810 6.070 13.980 6.240 ;
        RECT 14.150 6.070 14.320 6.240 ;
        RECT 14.490 6.070 14.660 6.240 ;
        RECT 14.830 6.070 15.000 6.240 ;
        RECT 15.170 6.070 15.340 6.240 ;
        RECT 15.510 6.070 15.680 6.240 ;
        RECT 15.850 6.070 16.020 6.240 ;
        RECT 16.190 6.070 16.360 6.240 ;
        RECT 16.530 6.070 16.700 6.240 ;
        RECT 16.870 6.070 17.040 6.240 ;
        RECT 17.210 6.070 17.380 6.240 ;
        RECT 17.550 6.070 17.720 6.240 ;
        RECT 17.890 6.070 18.060 6.240 ;
        RECT 18.230 6.070 18.400 6.240 ;
        RECT 18.570 6.070 18.740 6.240 ;
        RECT 18.910 6.070 19.080 6.240 ;
        RECT 19.250 6.070 19.420 6.240 ;
        RECT 19.590 6.070 19.760 6.240 ;
        RECT 19.930 6.070 20.100 6.240 ;
        RECT 20.270 6.070 20.440 6.240 ;
        RECT 18.820 4.220 18.990 4.390 ;
        RECT 19.250 4.220 19.420 4.390 ;
      LAYER met1 ;
        RECT 0.000 5.920 20.660 6.400 ;
        RECT 18.760 4.460 19.460 5.920 ;
        RECT 18.760 4.160 19.480 4.460 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.600 1.170 3.150 1.680 ;
        RECT 0.600 0.320 3.900 1.170 ;
        RECT 10.550 1.150 11.390 1.600 ;
        RECT 10.550 0.310 12.410 1.150 ;
      LAYER li1 ;
        RECT 3.220 0.320 3.900 0.730 ;
        RECT 11.600 0.320 12.410 0.820 ;
        RECT 0.000 0.150 20.670 0.320 ;
      LAYER mcon ;
        RECT 0.210 0.150 0.380 0.320 ;
        RECT 0.550 0.150 0.720 0.320 ;
        RECT 0.890 0.150 1.060 0.320 ;
        RECT 1.230 0.150 1.400 0.320 ;
        RECT 1.570 0.150 1.740 0.320 ;
        RECT 1.910 0.150 2.080 0.320 ;
        RECT 2.250 0.150 2.420 0.320 ;
        RECT 2.590 0.150 2.760 0.320 ;
        RECT 2.930 0.150 3.100 0.320 ;
        RECT 3.270 0.150 3.440 0.320 ;
        RECT 3.610 0.150 3.780 0.320 ;
        RECT 3.950 0.150 4.120 0.320 ;
        RECT 4.290 0.150 4.460 0.320 ;
        RECT 4.630 0.150 4.800 0.320 ;
        RECT 4.970 0.150 5.140 0.320 ;
        RECT 5.310 0.150 5.480 0.320 ;
        RECT 5.650 0.150 5.820 0.320 ;
        RECT 5.990 0.150 6.160 0.320 ;
        RECT 6.330 0.150 6.500 0.320 ;
        RECT 6.670 0.150 6.840 0.320 ;
        RECT 7.010 0.150 7.180 0.320 ;
        RECT 7.350 0.150 7.520 0.320 ;
        RECT 7.690 0.150 7.860 0.320 ;
        RECT 8.030 0.150 8.200 0.320 ;
        RECT 8.370 0.150 8.540 0.320 ;
        RECT 8.710 0.150 8.880 0.320 ;
        RECT 9.050 0.150 9.220 0.320 ;
        RECT 9.390 0.150 9.560 0.320 ;
        RECT 9.730 0.150 9.900 0.320 ;
        RECT 10.070 0.150 10.240 0.320 ;
        RECT 10.410 0.150 10.580 0.320 ;
        RECT 10.750 0.150 10.920 0.320 ;
        RECT 11.090 0.150 11.260 0.320 ;
        RECT 11.430 0.150 11.600 0.320 ;
        RECT 11.770 0.150 11.940 0.320 ;
        RECT 12.110 0.150 12.280 0.320 ;
        RECT 12.450 0.150 12.620 0.320 ;
        RECT 12.790 0.150 12.960 0.320 ;
        RECT 13.130 0.150 13.300 0.320 ;
        RECT 13.470 0.150 13.640 0.320 ;
        RECT 13.810 0.150 13.980 0.320 ;
        RECT 14.150 0.150 14.320 0.320 ;
        RECT 14.490 0.150 14.660 0.320 ;
        RECT 14.830 0.150 15.000 0.320 ;
        RECT 15.170 0.150 15.340 0.320 ;
        RECT 15.510 0.150 15.680 0.320 ;
        RECT 15.850 0.150 16.020 0.320 ;
        RECT 16.190 0.150 16.360 0.320 ;
        RECT 16.530 0.150 16.700 0.320 ;
        RECT 16.870 0.150 17.040 0.320 ;
        RECT 17.210 0.150 17.380 0.320 ;
        RECT 17.550 0.150 17.720 0.320 ;
        RECT 17.890 0.150 18.060 0.320 ;
        RECT 18.230 0.150 18.400 0.320 ;
        RECT 18.570 0.150 18.740 0.320 ;
        RECT 18.910 0.150 19.080 0.320 ;
        RECT 19.250 0.150 19.420 0.320 ;
        RECT 19.590 0.150 19.760 0.320 ;
        RECT 19.930 0.150 20.100 0.320 ;
      LAYER met1 ;
        RECT 0.000 0.000 20.670 0.480 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 1.300 3.270 6.370 3.550 ;
        RECT 8.600 3.270 9.020 3.520 ;
        RECT 0.010 3.100 10.410 3.270 ;
        RECT 11.140 3.100 20.660 3.270 ;
        RECT 0.930 2.040 1.120 3.100 ;
        RECT 2.170 2.040 2.360 3.100 ;
        RECT 4.010 2.730 9.250 3.100 ;
        RECT 12.080 2.820 19.570 3.100 ;
        RECT 4.010 2.720 9.420 2.730 ;
        RECT 3.880 2.550 9.420 2.720 ;
        RECT 4.620 2.540 9.420 2.550 ;
      LAYER mcon ;
        RECT 0.210 3.100 0.380 3.270 ;
        RECT 0.550 3.100 0.720 3.270 ;
        RECT 0.890 3.100 1.060 3.270 ;
        RECT 1.230 3.100 1.400 3.270 ;
        RECT 1.570 3.100 1.740 3.270 ;
        RECT 1.910 3.100 2.080 3.270 ;
        RECT 2.250 3.100 2.420 3.270 ;
        RECT 2.590 3.100 2.760 3.270 ;
        RECT 2.930 3.100 3.100 3.270 ;
        RECT 3.270 3.100 3.440 3.270 ;
        RECT 3.610 3.100 3.780 3.270 ;
        RECT 3.950 3.100 4.120 3.270 ;
        RECT 4.290 3.100 4.460 3.270 ;
        RECT 4.630 3.100 4.800 3.270 ;
        RECT 4.970 3.100 5.140 3.270 ;
        RECT 5.310 3.100 5.480 3.270 ;
        RECT 5.650 3.100 5.820 3.270 ;
        RECT 5.990 3.100 6.160 3.270 ;
        RECT 6.330 3.100 6.500 3.270 ;
        RECT 6.670 3.100 6.840 3.270 ;
        RECT 7.010 3.100 7.180 3.270 ;
        RECT 7.350 3.100 7.520 3.270 ;
        RECT 7.690 3.100 7.860 3.270 ;
        RECT 8.030 3.100 8.200 3.270 ;
        RECT 8.370 3.100 8.540 3.270 ;
        RECT 8.710 3.100 8.880 3.270 ;
        RECT 9.050 3.100 9.220 3.270 ;
        RECT 9.390 3.100 9.560 3.270 ;
        RECT 9.730 3.100 9.900 3.270 ;
        RECT 10.070 3.100 10.240 3.270 ;
        RECT 11.430 3.100 11.600 3.270 ;
        RECT 11.770 3.100 11.940 3.270 ;
        RECT 12.110 3.100 12.280 3.270 ;
        RECT 12.450 3.100 12.620 3.270 ;
        RECT 12.790 3.100 12.960 3.270 ;
        RECT 13.130 3.100 13.300 3.270 ;
        RECT 13.470 3.100 13.640 3.270 ;
        RECT 13.810 3.100 13.980 3.270 ;
        RECT 14.150 3.100 14.320 3.270 ;
        RECT 14.490 3.100 14.660 3.270 ;
        RECT 14.830 3.100 15.000 3.270 ;
        RECT 15.170 3.100 15.340 3.270 ;
        RECT 15.510 3.100 15.680 3.270 ;
        RECT 15.850 3.100 16.020 3.270 ;
        RECT 16.190 3.100 16.360 3.270 ;
        RECT 16.530 3.100 16.700 3.270 ;
        RECT 16.870 3.100 17.040 3.270 ;
        RECT 17.210 3.100 17.380 3.270 ;
        RECT 17.550 3.100 17.720 3.270 ;
        RECT 17.890 3.100 18.060 3.270 ;
        RECT 18.230 3.100 18.400 3.270 ;
        RECT 18.570 3.100 18.740 3.270 ;
        RECT 18.910 3.100 19.080 3.270 ;
        RECT 19.250 3.100 19.420 3.270 ;
        RECT 19.590 3.100 19.760 3.270 ;
        RECT 19.930 3.100 20.100 3.270 ;
      LAYER met1 ;
        RECT 0.010 2.960 20.660 3.440 ;
    END
  END GND
  PIN Up
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.225000 ;
    PORT
      LAYER li1 ;
        RECT 10.100 2.490 10.270 2.820 ;
        RECT 1.940 1.660 2.270 1.830 ;
      LAYER mcon ;
        RECT 10.100 2.570 10.270 2.740 ;
        RECT 2.020 1.660 2.190 1.830 ;
      LAYER met1 ;
        RECT 10.020 2.490 10.340 2.810 ;
        RECT 1.940 1.580 2.260 1.900 ;
      LAYER via ;
        RECT 10.050 2.520 10.310 2.780 ;
        RECT 1.970 1.610 2.230 1.870 ;
      LAYER met2 ;
        RECT 9.470 2.490 10.340 2.810 ;
        RECT 1.760 1.610 2.260 1.900 ;
        RECT 1.760 1.100 2.090 1.610 ;
        RECT 9.470 1.100 9.840 2.490 ;
        RECT 1.760 1.090 9.840 1.100 ;
        RECT 0.010 0.730 9.840 1.090 ;
    END
  END Up
  PIN Down
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.972000 ;
    PORT
      LAYER li1 ;
        RECT 2.040 4.030 2.210 4.360 ;
        RECT 0.700 1.660 1.030 1.830 ;
      LAYER mcon ;
        RECT 2.040 4.110 2.210 4.280 ;
        RECT 0.780 1.660 0.950 1.830 ;
      LAYER met1 ;
        RECT 1.960 4.030 2.280 4.350 ;
        RECT 0.710 1.580 1.030 1.900 ;
      LAYER via ;
        RECT 1.990 4.060 2.250 4.320 ;
        RECT 0.740 1.610 1.000 1.870 ;
      LAYER met2 ;
        RECT 1.840 4.330 2.280 4.350 ;
        RECT 0.600 4.030 2.280 4.330 ;
        RECT 0.600 3.970 2.270 4.030 ;
        RECT 0.600 2.720 0.920 3.970 ;
        RECT 0.010 2.410 0.920 2.720 ;
        RECT 0.600 1.900 0.920 2.410 ;
        RECT 0.600 1.580 1.030 1.900 ;
    END
  END Down
  PIN Out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.277200 ;
    PORT
      LAYER li1 ;
        RECT 11.850 3.870 20.660 4.020 ;
        RECT 10.610 3.490 20.660 3.870 ;
        RECT 10.610 3.480 11.960 3.490 ;
        RECT 10.610 2.730 10.960 3.480 ;
        RECT 10.540 2.560 10.960 2.730 ;
    END
  END Out
  PIN ENb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.700000 ;
    PORT
      LAYER li1 ;
        RECT 0.510 4.810 0.960 5.050 ;
    END
  END ENb
  OBS
      LAYER li1 ;
        RECT 1.720 5.390 20.480 5.580 ;
        RECT 8.370 5.340 8.750 5.390 ;
        RECT 9.630 5.340 10.010 5.390 ;
        RECT 11.870 5.340 12.250 5.390 ;
        RECT 1.220 4.900 2.160 5.090 ;
        RECT 2.480 4.900 20.480 5.090 ;
        RECT 8.370 4.850 8.750 4.900 ;
        RECT 9.630 4.850 10.010 4.900 ;
        RECT 2.480 4.350 9.020 4.520 ;
        RECT 11.870 4.500 12.250 4.900 ;
        RECT 7.990 3.760 8.240 4.350 ;
        RECT 8.430 4.300 9.020 4.350 ;
        RECT 11.850 4.310 12.270 4.500 ;
        RECT 8.480 4.250 9.020 4.300 ;
        RECT 8.550 4.190 9.020 4.250 ;
        RECT 8.600 3.830 9.020 4.190 ;
        RECT 11.220 4.080 11.550 4.250 ;
        RECT 7.950 3.590 8.280 3.760 ;
        RECT 1.410 2.500 1.670 2.760 ;
        RECT 0.930 0.690 1.120 1.450 ;
        RECT 1.410 0.730 1.600 2.500 ;
        RECT 2.650 1.740 2.840 2.400 ;
        RECT 3.370 2.060 4.320 2.250 ;
        RECT 10.540 2.220 10.960 2.250 ;
        RECT 9.990 2.170 10.960 2.220 ;
        RECT 4.620 1.980 10.960 2.170 ;
        RECT 2.170 0.700 2.360 1.460 ;
        RECT 2.650 1.380 4.310 1.740 ;
        RECT 4.620 1.500 11.150 1.690 ;
        RECT 2.650 0.740 2.840 1.380 ;
        RECT 10.170 1.100 10.420 1.500 ;
        RECT 10.600 1.460 11.150 1.500 ;
        RECT 10.670 1.420 11.150 1.460 ;
        RECT 10.720 1.370 11.150 1.420 ;
        RECT 10.730 1.170 11.150 1.370 ;
        RECT 10.130 0.930 10.460 1.100 ;
        RECT 10.730 0.690 11.150 0.900 ;
      LAYER mcon ;
        RECT 12.810 5.400 12.980 5.570 ;
        RECT 13.150 5.400 13.320 5.570 ;
        RECT 11.300 4.080 11.470 4.250 ;
        RECT 1.460 2.540 1.630 2.710 ;
        RECT 0.940 1.110 1.110 1.280 ;
        RECT 0.940 0.770 1.110 0.940 ;
        RECT 2.180 1.120 2.350 1.290 ;
        RECT 2.180 0.780 2.350 0.950 ;
        RECT 10.860 0.720 11.030 0.890 ;
      LAYER met1 ;
        RECT 12.750 5.340 13.430 5.630 ;
        RECT 11.220 4.020 11.540 4.320 ;
        RECT 1.380 2.460 1.700 2.780 ;
        RECT 12.680 1.540 13.470 2.290 ;
        RECT 0.900 0.990 1.150 1.340 ;
        RECT 2.140 0.990 2.390 1.350 ;
        RECT 12.680 0.990 13.160 1.540 ;
        RECT 0.900 0.690 13.160 0.990 ;
      LAYER via ;
        RECT 12.930 5.340 13.190 5.600 ;
        RECT 11.250 4.030 11.510 4.290 ;
        RECT 1.410 2.490 1.670 2.750 ;
        RECT 12.810 1.740 13.350 2.100 ;
      LAYER met2 ;
        RECT 8.700 4.000 11.540 4.320 ;
        RECT 8.700 3.000 9.170 4.000 ;
        RECT 1.380 2.600 9.170 3.000 ;
        RECT 1.380 2.460 1.700 2.600 ;
        RECT 12.780 1.710 13.390 5.630 ;
  END
END CP
END LIBRARY

