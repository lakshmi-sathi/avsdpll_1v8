magic
tech sky130A
timestamp 1605333160
<< nwell >>
rect -145 1311 381 1359
rect -145 1195 397 1311
rect -144 1188 397 1195
rect -144 1089 170 1188
rect 3 919 170 1089
rect -144 723 170 919
rect 3 658 170 723
rect 3 604 169 658
<< nmos >>
rect -82 1018 -67 1054
rect 246 1083 261 1125
rect -82 652 -67 688
rect 53 484 68 526
rect 190 496 205 537
rect 247 496 262 1036
rect 296 496 311 1036
<< pmos >>
rect -82 1114 -67 1186
rect -82 748 -67 820
rect 55 726 70 1266
rect 103 726 118 1266
rect 160 1224 175 1266
rect 317 1223 332 1265
rect 103 634 118 676
<< ndiff >>
rect -115 1045 -82 1054
rect -115 1028 -107 1045
rect -90 1028 -82 1045
rect -115 1018 -82 1028
rect -67 1045 -34 1054
rect -67 1028 -59 1045
rect -42 1028 -34 1045
rect -67 1018 -34 1028
rect 213 1113 246 1125
rect 213 1096 221 1113
rect 238 1096 246 1113
rect 213 1083 246 1096
rect 261 1113 294 1125
rect 261 1096 269 1113
rect 286 1096 294 1113
rect 261 1083 294 1096
rect 213 1029 247 1036
rect 213 1012 221 1029
rect 238 1012 247 1029
rect 213 995 247 1012
rect 213 978 221 995
rect 238 978 247 995
rect 213 961 247 978
rect 213 944 221 961
rect 238 944 247 961
rect 213 927 247 944
rect 213 910 221 927
rect 238 910 247 927
rect 213 893 247 910
rect 213 876 221 893
rect 238 876 247 893
rect 213 859 247 876
rect 213 842 221 859
rect 238 842 247 859
rect 213 825 247 842
rect 213 808 221 825
rect 238 808 247 825
rect 213 791 247 808
rect 213 774 221 791
rect 238 774 247 791
rect 213 757 247 774
rect 213 740 221 757
rect 238 740 247 757
rect 213 723 247 740
rect 213 706 221 723
rect 238 706 247 723
rect -115 679 -82 688
rect -115 662 -107 679
rect -90 662 -82 679
rect -115 652 -82 662
rect -67 679 -34 688
rect -67 662 -59 679
rect -42 662 -34 679
rect -67 652 -34 662
rect 213 689 247 706
rect 213 672 221 689
rect 238 672 247 689
rect 213 655 247 672
rect 213 638 221 655
rect 238 638 247 655
rect 213 621 247 638
rect 213 604 221 621
rect 238 604 247 621
rect 213 587 247 604
rect 213 570 221 587
rect 238 570 247 587
rect 213 553 247 570
rect 213 537 221 553
rect 20 514 53 526
rect 20 497 28 514
rect 45 497 53 514
rect 20 484 53 497
rect 68 515 101 526
rect 68 497 76 515
rect 93 497 101 515
rect 68 484 101 497
rect 157 525 190 537
rect 157 508 165 525
rect 182 508 190 525
rect 157 496 190 508
rect 205 536 221 537
rect 238 536 247 553
rect 205 519 247 536
rect 205 502 221 519
rect 238 502 247 519
rect 205 496 247 502
rect 262 1029 296 1036
rect 262 1012 270 1029
rect 287 1012 296 1029
rect 262 995 296 1012
rect 262 978 270 995
rect 287 978 296 995
rect 262 961 296 978
rect 262 944 270 961
rect 287 944 296 961
rect 262 927 296 944
rect 262 910 270 927
rect 287 910 296 927
rect 262 893 296 910
rect 262 876 270 893
rect 287 876 296 893
rect 262 859 296 876
rect 262 842 270 859
rect 287 842 296 859
rect 262 825 296 842
rect 262 808 270 825
rect 287 808 296 825
rect 262 791 296 808
rect 262 774 270 791
rect 287 774 296 791
rect 262 757 296 774
rect 262 740 270 757
rect 287 740 296 757
rect 262 723 296 740
rect 262 706 270 723
rect 287 706 296 723
rect 262 689 296 706
rect 262 672 270 689
rect 287 672 296 689
rect 262 655 296 672
rect 262 638 270 655
rect 287 638 296 655
rect 262 621 296 638
rect 262 604 270 621
rect 287 604 296 621
rect 262 587 296 604
rect 262 570 270 587
rect 287 570 296 587
rect 262 553 296 570
rect 262 536 270 553
rect 287 536 296 553
rect 262 519 296 536
rect 262 502 270 519
rect 287 502 296 519
rect 262 496 296 502
rect 311 1029 344 1036
rect 311 1012 319 1029
rect 336 1012 344 1029
rect 311 995 344 1012
rect 311 978 319 995
rect 336 978 344 995
rect 311 961 344 978
rect 311 944 319 961
rect 336 944 344 961
rect 311 927 344 944
rect 311 910 319 927
rect 336 910 344 927
rect 311 893 344 910
rect 311 876 319 893
rect 336 876 344 893
rect 311 859 344 876
rect 311 842 319 859
rect 336 842 344 859
rect 311 825 344 842
rect 311 808 319 825
rect 336 808 344 825
rect 311 791 344 808
rect 311 774 319 791
rect 336 774 344 791
rect 311 757 344 774
rect 311 740 319 757
rect 336 740 344 757
rect 311 723 344 740
rect 311 706 319 723
rect 336 706 344 723
rect 311 689 344 706
rect 311 672 319 689
rect 336 672 344 689
rect 311 655 344 672
rect 311 638 319 655
rect 336 638 344 655
rect 311 621 344 638
rect 311 604 319 621
rect 336 604 344 621
rect 311 587 344 604
rect 311 570 319 587
rect 336 570 344 587
rect 311 553 344 570
rect 311 536 319 553
rect 336 536 344 553
rect 311 519 344 536
rect 311 502 319 519
rect 336 502 344 519
rect 311 496 344 502
<< pdiff >>
rect 22 1258 55 1266
rect 22 1241 30 1258
rect 47 1241 55 1258
rect 22 1224 55 1241
rect 22 1207 30 1224
rect 47 1207 55 1224
rect 22 1190 55 1207
rect -116 1182 -82 1186
rect -116 1165 -107 1182
rect -90 1165 -82 1182
rect -116 1148 -82 1165
rect -116 1131 -107 1148
rect -90 1131 -82 1148
rect -116 1114 -82 1131
rect -67 1169 -35 1186
rect -67 1152 -59 1169
rect -42 1152 -35 1169
rect -67 1135 -35 1152
rect -67 1118 -59 1135
rect -42 1118 -35 1135
rect -67 1114 -35 1118
rect 22 1173 30 1190
rect 47 1173 55 1190
rect 22 1156 55 1173
rect 22 1139 30 1156
rect 47 1139 55 1156
rect 22 1122 55 1139
rect 22 1105 30 1122
rect 47 1105 55 1122
rect 22 1088 55 1105
rect 22 1071 30 1088
rect 47 1071 55 1088
rect 22 1054 55 1071
rect 22 1037 30 1054
rect 47 1037 55 1054
rect 22 1020 55 1037
rect 22 1003 30 1020
rect 47 1003 55 1020
rect 22 986 55 1003
rect 22 969 30 986
rect 47 969 55 986
rect 22 952 55 969
rect 22 935 30 952
rect 47 935 55 952
rect 22 918 55 935
rect 22 901 30 918
rect 47 901 55 918
rect 22 884 55 901
rect 22 867 30 884
rect 47 867 55 884
rect 22 850 55 867
rect 22 833 30 850
rect 47 833 55 850
rect -116 816 -82 820
rect -116 799 -107 816
rect -90 799 -82 816
rect -116 782 -82 799
rect -116 765 -107 782
rect -90 765 -82 782
rect -116 748 -82 765
rect -67 803 -35 820
rect -67 786 -59 803
rect -42 786 -35 803
rect -67 769 -35 786
rect -67 752 -59 769
rect -42 752 -35 769
rect -67 748 -35 752
rect 22 816 55 833
rect 22 799 30 816
rect 47 799 55 816
rect 22 782 55 799
rect 22 765 30 782
rect 47 765 55 782
rect 22 748 55 765
rect 22 731 30 748
rect 47 731 55 748
rect 22 726 55 731
rect 70 1258 103 1266
rect 70 1241 78 1258
rect 95 1241 103 1258
rect 70 1224 103 1241
rect 70 1207 78 1224
rect 95 1207 103 1224
rect 70 1190 103 1207
rect 70 1173 78 1190
rect 95 1173 103 1190
rect 70 1156 103 1173
rect 70 1139 78 1156
rect 95 1139 103 1156
rect 70 1122 103 1139
rect 70 1105 78 1122
rect 95 1105 103 1122
rect 70 1088 103 1105
rect 70 1071 78 1088
rect 95 1071 103 1088
rect 70 1054 103 1071
rect 70 1037 78 1054
rect 95 1037 103 1054
rect 70 1020 103 1037
rect 70 1003 78 1020
rect 95 1003 103 1020
rect 70 986 103 1003
rect 70 969 78 986
rect 95 969 103 986
rect 70 952 103 969
rect 70 935 78 952
rect 95 935 103 952
rect 70 918 103 935
rect 70 901 78 918
rect 95 901 103 918
rect 70 884 103 901
rect 70 867 78 884
rect 95 867 103 884
rect 70 850 103 867
rect 70 833 78 850
rect 95 833 103 850
rect 70 816 103 833
rect 70 799 78 816
rect 95 799 103 816
rect 70 782 103 799
rect 70 765 78 782
rect 95 765 103 782
rect 70 748 103 765
rect 70 731 78 748
rect 95 731 103 748
rect 70 726 103 731
rect 118 1258 160 1266
rect 118 1241 126 1258
rect 143 1241 160 1258
rect 118 1224 160 1241
rect 175 1254 208 1266
rect 175 1237 183 1254
rect 200 1237 208 1254
rect 175 1224 208 1237
rect 284 1253 317 1265
rect 284 1236 292 1253
rect 309 1236 317 1253
rect 118 1207 126 1224
rect 143 1207 152 1224
rect 284 1223 317 1236
rect 332 1253 366 1265
rect 332 1236 340 1253
rect 357 1236 366 1253
rect 332 1223 366 1236
rect 118 1190 152 1207
rect 118 1173 126 1190
rect 143 1173 152 1190
rect 118 1156 152 1173
rect 118 1139 126 1156
rect 143 1139 152 1156
rect 118 1122 152 1139
rect 118 1105 126 1122
rect 143 1105 152 1122
rect 118 1088 152 1105
rect 118 1071 126 1088
rect 143 1071 152 1088
rect 118 1054 152 1071
rect 118 1037 126 1054
rect 143 1037 152 1054
rect 118 1020 152 1037
rect 118 1003 126 1020
rect 143 1003 152 1020
rect 118 986 152 1003
rect 118 969 126 986
rect 143 969 152 986
rect 118 952 152 969
rect 118 935 126 952
rect 143 935 152 952
rect 118 918 152 935
rect 118 901 126 918
rect 143 901 152 918
rect 118 884 152 901
rect 118 867 126 884
rect 143 867 152 884
rect 118 850 152 867
rect 118 833 126 850
rect 143 833 152 850
rect 118 816 152 833
rect 118 799 126 816
rect 143 799 152 816
rect 118 782 152 799
rect 118 765 126 782
rect 143 765 152 782
rect 118 748 152 765
rect 118 731 126 748
rect 143 731 152 748
rect 118 726 152 731
rect 70 664 103 676
rect 70 647 78 664
rect 95 647 103 664
rect 70 634 103 647
rect 118 664 151 676
rect 118 647 126 664
rect 143 647 151 664
rect 118 634 151 647
<< ndiffc >>
rect -107 1028 -90 1045
rect -59 1028 -42 1045
rect 221 1096 238 1113
rect 269 1096 286 1113
rect 221 1012 238 1029
rect 221 978 238 995
rect 221 944 238 961
rect 221 910 238 927
rect 221 876 238 893
rect 221 842 238 859
rect 221 808 238 825
rect 221 774 238 791
rect 221 740 238 757
rect 221 706 238 723
rect -107 662 -90 679
rect -59 662 -42 679
rect 221 672 238 689
rect 221 638 238 655
rect 221 604 238 621
rect 221 570 238 587
rect 28 497 45 514
rect 76 497 93 515
rect 165 508 182 525
rect 221 536 238 553
rect 221 502 238 519
rect 270 1012 287 1029
rect 270 978 287 995
rect 270 944 287 961
rect 270 910 287 927
rect 270 876 287 893
rect 270 842 287 859
rect 270 808 287 825
rect 270 774 287 791
rect 270 740 287 757
rect 270 706 287 723
rect 270 672 287 689
rect 270 638 287 655
rect 270 604 287 621
rect 270 570 287 587
rect 270 536 287 553
rect 270 502 287 519
rect 319 1012 336 1029
rect 319 978 336 995
rect 319 944 336 961
rect 319 910 336 927
rect 319 876 336 893
rect 319 842 336 859
rect 319 808 336 825
rect 319 774 336 791
rect 319 740 336 757
rect 319 706 336 723
rect 319 672 336 689
rect 319 638 336 655
rect 319 604 336 621
rect 319 570 336 587
rect 319 536 336 553
rect 319 502 336 519
<< pdiffc >>
rect 30 1241 47 1258
rect 30 1207 47 1224
rect -107 1165 -90 1182
rect -107 1131 -90 1148
rect -59 1152 -42 1169
rect -59 1118 -42 1135
rect 30 1173 47 1190
rect 30 1139 47 1156
rect 30 1105 47 1122
rect 30 1071 47 1088
rect 30 1037 47 1054
rect 30 1003 47 1020
rect 30 969 47 986
rect 30 935 47 952
rect 30 901 47 918
rect 30 867 47 884
rect 30 833 47 850
rect -107 799 -90 816
rect -107 765 -90 782
rect -59 786 -42 803
rect -59 752 -42 769
rect 30 799 47 816
rect 30 765 47 782
rect 30 731 47 748
rect 78 1241 95 1258
rect 78 1207 95 1224
rect 78 1173 95 1190
rect 78 1139 95 1156
rect 78 1105 95 1122
rect 78 1071 95 1088
rect 78 1037 95 1054
rect 78 1003 95 1020
rect 78 969 95 986
rect 78 935 95 952
rect 78 901 95 918
rect 78 867 95 884
rect 78 833 95 850
rect 78 799 95 816
rect 78 765 95 782
rect 78 731 95 748
rect 126 1241 143 1258
rect 183 1237 200 1254
rect 292 1236 309 1253
rect 126 1207 143 1224
rect 340 1236 357 1253
rect 126 1173 143 1190
rect 126 1139 143 1156
rect 126 1105 143 1122
rect 126 1071 143 1088
rect 126 1037 143 1054
rect 126 1003 143 1020
rect 126 969 143 986
rect 126 935 143 952
rect 126 901 143 918
rect 126 867 143 884
rect 126 833 143 850
rect 126 799 143 816
rect 126 765 143 782
rect 126 731 143 748
rect 78 647 95 664
rect 126 647 143 664
<< psubdiff >>
rect -121 972 -109 990
rect -92 972 -80 990
rect -121 606 -109 624
rect -92 606 -80 624
rect -124 415 -112 432
rect -95 415 -83 432
rect -42 415 -30 432
rect -13 415 -1 432
rect 40 415 52 432
rect 69 415 81 432
rect 122 415 134 432
rect 151 415 163 432
rect 204 415 216 432
rect 233 415 245 432
rect 286 415 298 432
rect 315 415 327 432
<< nsubdiff >>
rect -117 1324 -105 1341
rect -88 1324 -75 1341
rect -33 1324 -21 1341
rect -4 1324 9 1341
rect 51 1324 63 1341
rect 80 1324 93 1341
rect 135 1324 147 1341
rect 164 1324 177 1341
rect 219 1324 231 1341
rect 248 1324 261 1341
rect 303 1324 315 1341
rect 332 1324 345 1341
rect -119 1218 -107 1235
rect -90 1218 -78 1235
rect -119 852 -107 869
rect -90 852 -78 869
<< psubdiffcont >>
rect -109 972 -92 990
rect -109 606 -92 624
rect -112 415 -95 432
rect -30 415 -13 432
rect 52 415 69 432
rect 134 415 151 432
rect 216 415 233 432
rect 298 415 315 432
<< nsubdiffcont >>
rect -105 1324 -88 1341
rect -21 1324 -4 1341
rect 63 1324 80 1341
rect 147 1324 164 1341
rect 231 1324 248 1341
rect 315 1324 332 1341
rect -107 1218 -90 1235
rect -107 852 -90 869
<< poly >>
rect 103 1279 241 1296
rect 55 1266 70 1279
rect 103 1266 118 1279
rect 160 1278 241 1279
rect 160 1266 175 1278
rect -82 1186 -67 1199
rect -82 1100 -67 1114
rect -111 1090 -67 1100
rect -111 1073 -103 1090
rect -86 1073 -67 1090
rect -111 1067 -67 1073
rect -82 1054 -67 1067
rect -82 1004 -67 1018
rect -82 820 -67 833
rect -82 733 -67 748
rect -116 724 -67 733
rect 222 1263 241 1278
rect 317 1265 332 1278
rect 222 1253 251 1263
rect 222 1236 228 1253
rect 245 1236 251 1253
rect 222 1224 251 1236
rect 160 1211 175 1224
rect 317 1210 332 1223
rect 317 1203 392 1210
rect 317 1194 367 1203
rect 359 1186 367 1194
rect 384 1186 392 1203
rect 359 1181 392 1186
rect 237 1162 272 1168
rect 237 1145 246 1162
rect 263 1145 272 1162
rect 237 1140 272 1145
rect 246 1125 261 1140
rect 246 1070 261 1083
rect 247 1036 262 1049
rect 296 1036 311 1049
rect -116 707 -106 724
rect -89 707 -67 724
rect 55 714 70 726
rect -116 702 -67 707
rect -82 688 -67 702
rect -7 694 70 714
rect 103 713 118 726
rect -82 638 -67 652
rect -7 636 15 694
rect 103 676 118 690
rect -29 625 15 636
rect -29 601 -24 625
rect -1 601 15 625
rect 103 621 118 634
rect 103 608 179 621
rect 103 606 157 608
rect -29 592 15 601
rect 152 591 157 606
rect 174 591 179 608
rect 152 586 179 591
rect 157 583 174 586
rect 36 569 69 575
rect 36 552 44 569
rect 61 552 69 569
rect 36 547 69 552
rect 53 526 68 547
rect 115 531 142 542
rect 190 537 205 550
rect 115 514 120 531
rect 137 514 142 531
rect 115 506 142 514
rect 122 486 142 506
rect 369 533 396 541
rect 369 516 374 533
rect 391 516 396 533
rect 369 508 396 516
rect 190 486 205 496
rect 247 486 262 496
rect 53 471 68 484
rect 122 471 262 486
rect 296 486 311 496
rect 369 486 386 508
rect 296 471 386 486
<< polycont >>
rect -103 1073 -86 1090
rect 228 1236 245 1253
rect 367 1186 384 1203
rect 246 1145 263 1162
rect -106 707 -89 724
rect -24 601 -1 625
rect 157 591 174 608
rect 44 552 61 569
rect 120 514 137 531
rect 374 516 391 533
<< locali >>
rect -154 1341 423 1361
rect -154 1324 -105 1341
rect -88 1324 -21 1341
rect -4 1324 63 1341
rect 80 1324 147 1341
rect 164 1324 231 1341
rect 248 1324 315 1341
rect 332 1324 423 1341
rect -154 1311 423 1324
rect 29 1258 48 1266
rect -108 1235 -89 1247
rect -108 1218 -107 1235
rect -90 1218 -89 1235
rect -108 1182 -89 1218
rect 29 1241 30 1258
rect 47 1241 48 1258
rect 29 1224 48 1241
rect 29 1207 30 1224
rect 47 1207 48 1224
rect 29 1190 48 1207
rect -108 1165 -107 1182
rect -90 1165 -89 1182
rect -108 1148 -89 1165
rect -108 1131 -107 1148
rect -90 1131 -89 1148
rect -108 1114 -89 1131
rect -60 1169 -41 1186
rect -60 1152 -59 1169
rect -42 1152 -41 1169
rect -60 1135 -41 1152
rect -60 1118 -59 1135
rect -42 1118 -41 1135
rect -60 1094 -41 1118
rect 29 1173 30 1190
rect 47 1173 48 1190
rect 29 1156 48 1173
rect 29 1139 30 1156
rect 47 1139 48 1156
rect 29 1122 48 1139
rect 29 1105 30 1122
rect 47 1105 48 1122
rect -152 1090 -78 1093
rect -152 1073 -103 1090
rect -86 1073 -78 1090
rect -152 1071 -78 1073
rect -60 1090 -8 1094
rect -60 1073 -32 1090
rect -15 1073 -8 1090
rect -151 944 -131 1071
rect -60 1068 -8 1073
rect 29 1088 48 1105
rect 29 1071 30 1088
rect 47 1071 48 1088
rect -108 1045 -89 1054
rect -108 1028 -107 1045
rect -90 1028 -89 1045
rect -108 1018 -89 1028
rect -60 1045 -41 1068
rect -60 1028 -59 1045
rect -42 1028 -41 1045
rect -60 1018 -41 1028
rect 29 1054 48 1071
rect 29 1037 30 1054
rect 47 1037 48 1054
rect 29 1020 48 1037
rect -108 1007 -90 1018
rect -110 990 -90 1007
rect -110 972 -109 990
rect -92 972 -90 990
rect -110 964 -90 972
rect 29 1003 30 1020
rect 47 1003 48 1020
rect 29 986 48 1003
rect 29 969 30 986
rect 47 969 48 986
rect 29 952 48 969
rect -151 938 10 944
rect -151 907 11 938
rect -108 869 -89 881
rect -108 852 -107 869
rect -90 852 -89 869
rect -108 816 -89 852
rect -14 843 11 907
rect 29 935 30 952
rect 47 935 48 952
rect 29 918 48 935
rect 29 901 30 918
rect 47 901 48 918
rect 29 884 48 901
rect 29 867 30 884
rect 47 867 48 884
rect 29 850 48 867
rect -108 799 -107 816
rect -90 799 -89 816
rect -108 782 -89 799
rect -108 765 -107 782
rect -90 765 -89 782
rect -108 748 -89 765
rect -60 803 -41 820
rect -60 786 -59 803
rect -42 786 -41 803
rect -60 769 -41 786
rect -60 752 -59 769
rect -42 752 -41 769
rect -60 727 -41 752
rect -114 707 -106 724
rect -89 707 -81 724
rect -108 679 -89 688
rect -108 662 -107 679
rect -90 662 -89 679
rect -108 652 -89 662
rect -60 679 -41 704
rect -60 662 -59 679
rect -42 662 -41 679
rect -60 652 -41 662
rect -108 641 -90 652
rect -110 624 -90 641
rect -14 636 10 843
rect -110 606 -109 624
rect -92 606 -90 624
rect -110 598 -90 606
rect -24 625 10 636
rect -1 601 10 625
rect -24 591 10 601
rect 29 833 30 850
rect 47 833 48 850
rect 29 816 48 833
rect 29 799 30 816
rect 47 799 48 816
rect 29 782 48 799
rect 29 765 30 782
rect 47 765 48 782
rect 29 748 48 765
rect 29 731 30 748
rect 47 731 48 748
rect 29 588 48 731
rect 77 1258 96 1266
rect 77 1241 78 1258
rect 95 1241 96 1258
rect 77 1224 96 1241
rect 77 1207 78 1224
rect 95 1207 96 1224
rect 77 1190 96 1207
rect 77 1173 78 1190
rect 95 1173 96 1190
rect 77 1156 96 1173
rect 77 1139 78 1156
rect 95 1139 96 1156
rect 77 1122 96 1139
rect 77 1105 78 1122
rect 95 1105 96 1122
rect 77 1088 96 1105
rect 77 1071 78 1088
rect 95 1071 96 1088
rect 77 1054 96 1071
rect 77 1037 78 1054
rect 95 1037 96 1054
rect 77 1020 96 1037
rect 77 1003 78 1020
rect 95 1003 96 1020
rect 77 986 96 1003
rect 77 969 78 986
rect 95 969 96 986
rect 77 952 96 969
rect 77 935 78 952
rect 95 935 96 952
rect 77 918 96 935
rect 77 901 78 918
rect 95 901 96 918
rect 77 884 96 901
rect 77 867 78 884
rect 95 867 96 884
rect 77 850 96 867
rect 77 833 78 850
rect 95 833 96 850
rect 77 816 96 833
rect 77 799 78 816
rect 95 799 96 816
rect 77 782 96 799
rect 77 765 78 782
rect 95 765 96 782
rect 77 748 96 765
rect 77 731 78 748
rect 95 731 96 748
rect 77 664 96 731
rect 125 1258 144 1311
rect 272 1302 330 1311
rect 281 1278 320 1302
rect 125 1241 126 1258
rect 143 1241 144 1258
rect 125 1224 144 1241
rect 183 1257 200 1266
rect 227 1257 246 1261
rect 183 1254 246 1257
rect 200 1253 246 1254
rect 200 1237 228 1253
rect 183 1236 228 1237
rect 245 1236 246 1253
rect 183 1235 246 1236
rect 183 1224 200 1235
rect 227 1226 246 1235
rect 291 1253 310 1278
rect 291 1236 292 1253
rect 309 1236 310 1253
rect 125 1207 126 1224
rect 143 1207 144 1224
rect 291 1223 310 1236
rect 339 1256 375 1265
rect 339 1253 385 1256
rect 339 1236 340 1253
rect 357 1236 385 1253
rect 339 1223 385 1236
rect 125 1190 144 1207
rect 125 1173 126 1190
rect 143 1173 144 1190
rect 125 1156 144 1173
rect 366 1203 385 1223
rect 366 1186 367 1203
rect 384 1186 385 1203
rect 125 1139 126 1156
rect 143 1139 144 1156
rect 238 1145 246 1162
rect 263 1145 272 1162
rect 366 1161 385 1186
rect 125 1122 144 1139
rect 318 1140 385 1161
rect 125 1105 126 1122
rect 143 1105 144 1122
rect 125 1088 144 1105
rect 125 1071 126 1088
rect 143 1071 144 1088
rect 220 1113 239 1125
rect 220 1096 221 1113
rect 238 1096 239 1113
rect 220 1083 239 1096
rect 268 1113 287 1125
rect 268 1096 269 1113
rect 286 1096 287 1113
rect 268 1083 287 1096
rect 125 1054 144 1071
rect 125 1037 126 1054
rect 143 1037 144 1054
rect 269 1037 287 1083
rect 125 1020 144 1037
rect 125 1003 126 1020
rect 143 1003 144 1020
rect 125 986 144 1003
rect 125 969 126 986
rect 143 969 144 986
rect 125 952 144 969
rect 125 935 126 952
rect 143 935 144 952
rect 125 918 144 935
rect 125 901 126 918
rect 143 901 144 918
rect 125 884 144 901
rect 125 867 126 884
rect 143 867 144 884
rect 125 850 144 867
rect 125 833 126 850
rect 143 833 144 850
rect 125 816 144 833
rect 125 799 126 816
rect 143 799 144 816
rect 125 782 144 799
rect 125 765 126 782
rect 143 765 144 782
rect 125 748 144 765
rect 125 731 126 748
rect 143 731 144 748
rect 125 723 144 731
rect 220 1029 239 1037
rect 220 1012 221 1029
rect 238 1012 239 1029
rect 220 995 239 1012
rect 220 978 221 995
rect 238 978 239 995
rect 220 961 239 978
rect 220 944 221 961
rect 238 944 239 961
rect 220 927 239 944
rect 220 910 221 927
rect 238 910 239 927
rect 220 893 239 910
rect 220 876 221 893
rect 238 876 239 893
rect 220 859 239 876
rect 220 842 221 859
rect 238 842 239 859
rect 220 825 239 842
rect 220 808 221 825
rect 238 808 239 825
rect 220 791 239 808
rect 220 774 221 791
rect 238 774 239 791
rect 220 757 239 774
rect 220 740 221 757
rect 238 740 239 757
rect 220 723 239 740
rect 220 706 221 723
rect 238 706 239 723
rect 220 689 239 706
rect 77 647 78 664
rect 95 647 96 664
rect 77 634 96 647
rect 125 664 144 676
rect 125 647 126 664
rect 143 647 144 664
rect 125 634 144 647
rect 220 672 221 689
rect 238 672 239 689
rect 220 655 239 672
rect 220 638 221 655
rect 238 638 239 655
rect 220 621 239 638
rect 157 608 174 616
rect 28 575 49 588
rect 157 583 174 591
rect 220 604 221 621
rect 238 604 239 621
rect 220 587 239 604
rect 28 570 64 575
rect 220 570 221 587
rect 238 570 239 587
rect 28 569 69 570
rect 28 555 44 569
rect 25 552 44 555
rect 61 552 69 569
rect 25 551 69 552
rect 220 553 239 570
rect 25 548 64 551
rect 22 547 64 548
rect 22 537 46 547
rect 20 514 46 537
rect 118 531 139 541
rect 20 497 28 514
rect 45 497 46 514
rect 20 484 46 497
rect 76 515 93 526
rect 118 514 120 531
rect 137 528 139 531
rect 164 528 183 537
rect 137 525 183 528
rect 137 514 165 525
rect 118 508 165 514
rect 182 508 183 525
rect 118 505 183 508
rect 76 481 93 497
rect 164 496 183 505
rect 220 536 221 553
rect 238 536 239 553
rect 220 519 239 536
rect 220 502 221 519
rect 238 502 239 519
rect 76 480 101 481
rect 65 473 101 480
rect 64 462 103 473
rect 64 461 109 462
rect 58 449 109 461
rect 220 449 239 502
rect 269 1029 288 1037
rect 269 1012 270 1029
rect 287 1012 288 1029
rect 269 995 288 1012
rect 269 978 270 995
rect 287 978 288 995
rect 269 961 288 978
rect 269 944 270 961
rect 287 944 288 961
rect 269 927 288 944
rect 269 910 270 927
rect 287 910 288 927
rect 269 893 288 910
rect 269 876 270 893
rect 287 876 288 893
rect 269 859 288 876
rect 269 842 270 859
rect 287 842 288 859
rect 269 825 288 842
rect 269 808 270 825
rect 287 808 288 825
rect 269 791 288 808
rect 269 774 270 791
rect 287 774 288 791
rect 269 757 288 774
rect 269 740 270 757
rect 287 740 288 757
rect 269 723 288 740
rect 269 706 270 723
rect 287 706 288 723
rect 269 689 288 706
rect 269 672 270 689
rect 287 672 288 689
rect 269 655 288 672
rect 269 638 270 655
rect 287 638 288 655
rect 269 621 288 638
rect 269 604 270 621
rect 287 604 288 621
rect 269 587 288 604
rect 269 570 270 587
rect 287 570 288 587
rect 269 553 288 570
rect 269 536 270 553
rect 287 536 288 553
rect 269 519 288 536
rect 269 502 270 519
rect 287 502 288 519
rect 269 494 288 502
rect 318 1029 337 1140
rect 318 1012 319 1029
rect 336 1012 337 1029
rect 318 995 337 1012
rect 318 978 319 995
rect 336 978 337 995
rect 318 961 337 978
rect 318 944 319 961
rect 336 944 337 961
rect 318 927 337 944
rect 318 910 319 927
rect 336 910 337 927
rect 318 893 337 910
rect 318 876 319 893
rect 336 876 337 893
rect 375 915 411 923
rect 375 887 376 915
rect 404 887 411 915
rect 375 878 411 887
rect 318 859 337 876
rect 318 842 319 859
rect 336 842 337 859
rect 318 825 337 842
rect 318 808 319 825
rect 336 808 337 825
rect 318 791 337 808
rect 318 774 319 791
rect 336 774 337 791
rect 318 757 337 774
rect 318 740 319 757
rect 336 740 337 757
rect 318 723 337 740
rect 318 706 319 723
rect 336 706 337 723
rect 318 689 337 706
rect 318 672 319 689
rect 336 672 337 689
rect 318 655 337 672
rect 318 638 319 655
rect 336 638 337 655
rect 318 621 337 638
rect 318 604 319 621
rect 336 604 337 621
rect 318 587 337 604
rect 318 570 319 587
rect 336 570 337 587
rect 318 553 337 570
rect 318 536 319 553
rect 336 536 337 553
rect 318 519 337 536
rect 318 502 319 519
rect 336 502 337 519
rect 374 533 391 541
rect 374 508 391 516
rect 318 494 337 502
rect -155 432 424 449
rect -155 415 -112 432
rect -95 415 -30 432
rect -13 415 52 432
rect 69 415 134 432
rect 151 415 216 432
rect 233 415 298 432
rect 315 415 424 432
rect -155 401 424 415
<< viali >>
rect -32 1073 -15 1090
rect -106 707 -89 724
rect -60 704 -39 727
rect 246 1145 263 1162
rect 221 1096 238 1113
rect 126 647 143 664
rect 157 591 174 608
rect 376 887 404 915
rect 374 516 391 533
<< metal1 >>
rect 61 1162 269 1168
rect 61 1145 246 1162
rect 263 1145 269 1162
rect 61 1139 269 1145
rect 61 1134 203 1139
rect -40 1095 -7 1098
rect -40 1069 -37 1095
rect -11 1069 -7 1095
rect -40 1066 -7 1069
rect 61 930 88 1134
rect 215 1113 409 1119
rect 215 1096 221 1113
rect 238 1096 409 1113
rect 215 1090 409 1096
rect -155 891 88 930
rect 372 915 409 1090
rect -155 824 -126 891
rect 372 887 376 915
rect 404 887 409 915
rect -155 731 -125 824
rect -155 724 -83 731
rect -155 707 -106 724
rect -89 707 -83 724
rect -155 702 -83 707
rect -67 727 -32 731
rect -67 704 -60 727
rect -39 704 -32 727
rect -67 549 -32 704
rect 372 670 409 887
rect 120 664 409 670
rect 120 647 126 664
rect 143 647 409 664
rect 120 641 409 647
rect 149 612 181 615
rect 149 586 152 612
rect 178 586 181 612
rect 149 583 181 586
rect -68 542 396 549
rect -68 533 397 542
rect -68 519 374 533
rect 368 516 374 519
rect 391 516 397 533
rect 368 510 397 516
<< via1 >>
rect -37 1090 -11 1095
rect -37 1073 -32 1090
rect -32 1073 -15 1090
rect -15 1073 -11 1090
rect -37 1069 -11 1073
rect 152 608 178 612
rect 152 591 157 608
rect 157 591 174 608
rect 174 591 178 608
rect 152 586 178 591
<< metal2 >>
rect -40 1095 -7 1098
rect -40 1069 -37 1095
rect -11 1069 179 1095
rect -40 1066 -7 1069
rect 152 615 179 1069
rect 149 612 181 615
rect 149 586 152 612
rect 178 586 181 612
rect 149 583 181 586
<< labels >>
rlabel locali -20 600 4 625 1 Down
port 1 n
rlabel metal1 376 886 404 916 1 Out
port 3 n
rlabel locali -154 1311 -154 1361 3 VDD
port 4 e
rlabel locali -155 401 -155 449 3 GND
port 5 e
rlabel metal1 -152 705 -128 729 1 Up
port 6 n
<< end >>
