*---------PLL---------
.include sky130nm.lib

xx1 clk_ref clk_vco_by_8 up down phase_detector
xx2 up down vin_vco charge_pump
xx3 vin_vco clk_out vcoscillator
c3 clk_vco_by_8 0 10f
xx5 clk_out 4 freqdiv2
xx6 4 3 freqdiv2
xx7 3 clk_vco_by_8 freqdiv2
*xm8 1 clk_out 6 1 sky130_fd_pr__pfet_01v8 l=150n w=720n 
*xm9 6 clk_out 0 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
*xm10 1 6 out 1 sky130_fd_pr__pfet_01v8 l=150n w=1440n 
*xm11 out 6 0 0 sky130_fd_pr__nfet_01v8 l=150n w=720n

v1 clk_ref 0 PULSE 0 1.8 10p 60p 60p 100ns 200ns
v2 1 0 1.8

*PD-----------------
.subckt phase_detector clk1 clk2 up down
xm1 1 clk1 3 1 sky130_fd_pr__pfet_01v8 l=150n w=420n 
xm2 3 clk1 4 0 sky130_fd_pr__nfet_01v8 l=150n w=420n
xm3 4 clk2 0 0 sky130_fd_pr__nfet_01v8 l=150n w=420n

xm4 1 clk2 6 1 sky130_fd_pr__pfet_01v8 l=150n w=420n 
xm5 6 clk2 7 0 sky130_fd_pr__nfet_01v8 l=150n w=420n
xm6 7 clk1 0 0 sky130_fd_pr__nfet_01v8 l=150n w=420n

xm7 8 clk1 3 0 sky130_fd_pr__nfet_01v8 l=150n w=1120n 
xm8 clk1 clk1 8 1 sky130_fd_pr__pfet_01v8 l=150n w=1120n

xm9 9 clk2 6 0 sky130_fd_pr__nfet_01v8 l=150n w=1120n
xm10 clk2 clk2 9 1 sky130_fd_pr__pfet_01v8 l=150n w=1120n

*buffer
xm11 1 8 10 1 sky130_fd_pr__pfet_01v8 l=150n w=720n 
xm12 10 8 0 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm15 1 10 up 1 sky130_fd_pr__pfet_01v8 l=150n w=720n 
xm16 up 10 0 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm13 1 9 11 1 sky130_fd_pr__pfet_01v8 l=150n w=720n 
xm17 11 9 0 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm18 1 11 down 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm14 down 11 0 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

*output cap
c1 8 0 0.35f
c2 9 0 0.35f

v1 1 0 1.8

.ends phase_detector
*--------------------

*CP-----------------
.subckt charge_pump up down out
xm1 upb up 0 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm2 downb down 0 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm3 1 down downb 1 sky130_fd_pr__pfet_01v8 l=150n w=1080n
xm4 1 up upb 1 sky130_fd_pr__pfet_01v8 l=150n w=1080n
xm5 upb 0 5 5 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm6 downb 0 4 4 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm7 3 4 3 3 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm8 0 1 1 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm9 out 1 3 3 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm10 3 down 0 0 sky130_fd_pr__nfet_01v8 l=150n w=30u
xm11 5 1 upb 5 sky130_fd_pr__pfet_01v8 l=150n w=1080n
xm12 4 1 downb 4 sky130_fd_pr__pfet_01v8 l=150n w=1080n
xm13 2 up 2 2 sky130_fd_pr__pfet_01v8 l=150n w=1080n
xm14 0 0 1 1 sky130_fd_pr__pfet_01v8 l=150n w=1080n
xm15 2 0 out 2 sky130_fd_pr__pfet_01v8 l=150n w=1080n
xm16 1 5 2 1 sky130_fd_pr__pfet_01v8 l=150n w=90u

*output cap
c1 out 0 1f

v1 1 0 1.8
.ends charge_pump
*--------------------

*LPF----------------
c1 vin_vco 0 200p
c2 5 0 500p
r1 vin_vco 5 500
*-------------------

*VCO----------------
.subckt vcoscillator vin vout
xm1 vp vn 0 0 sky130_fd_pr__nfet_01v8 l=200n w=400n
xm2 vp vp 1 1 sky130_fd_pr__pfet_01v8 l=200n w=2000n
r1 vn vin 1
*xu1 osc_fb Osc inv_20_10
xm3 1 osc_fb vout 1 sky130_fd_pr__pfet_01v8 l=150n w=2400n 
xm4 vout osc_fb 0 0 sky130_fd_pr__nfet_01v8 l=150n w=1200n
xx1 7 osc_fb vp vn cs_inv
xx2 6 7 vp vn cs_inv
xx3 5 6 vp vn cs_inv
xx4 4 5 vp vn cs_inv
xx5 3 4 vp vn cs_inv
xx6 2 3 vp vn cs_inv
xx7 osc_fb 2 vp vn cs_inv
*c1 vout 0 0.1f

v1 1 0 1.8
.ends vcoscillator

.subckt cs_inv in out vp vn
xm1 3 vn 0 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm2 2 vp 1 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm3 out in 2 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm4 out in 3 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

c1 out 0 1f
v1 1 0 1.8
.ends cs_inv
*----------------------

*FreqDiv by 2-----------
.subckt freqdiv2 clkin clkout 
xm1 1 5 2 1 sky130_fd_pr__pfet_01v8 l=150n w=3600n 
xm2 2 clkin 0 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm3 1 2 4 1 sky130_fd_pr__pfet_01v8 l=150n w=420n 
xm4 4 clkin 0 0 sky130_fd_pr__nfet_01v8 l=150n w=1120n

xm5 1 clkin 5 1 sky130_fd_pr__pfet_01v8 l=150n w=2400n 
xm6 5 4 0 0 sky130_fd_pr__nfet_01v8 l=150n w=4800n

*c1 5 0 0.1f

xm7 1 5 6 1 sky130_fd_pr__pfet_01v8 l=150n w=1120n 
xm8 6 5 0 0 sky130_fd_pr__nfet_01v8 l=150n w=560n

xm9 1 6 clkout 1 sky130_fd_pr__pfet_01v8 l=150n w=1120n 
xm10 clkout 6 0 0 sky130_fd_pr__nfet_01v8 l=150n w=560n


v1 1 0 1.8
.ends freqdiv2
*-----------------------


*simulation
.ic V(vin_vco) = 0
.control
tran 10ns 5us
*plot v(clk_ref)+8 v(up)+6 v(down)+4 v(vin_vco)+2 v(clk_out)
plot v(4)+2 v(clk_out) 

.endc
.end 