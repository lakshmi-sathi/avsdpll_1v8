magic
tech sky130A
timestamp 1607692587
<< nwell >>
rect 12 252 171 298
rect 12 144 346 252
<< pwell >>
rect 30 -15 71 4
<< nmos >>
rect 65 64 80 106
rect 171 64 186 106
rect 284 64 299 106
<< pmos >>
rect 65 162 80 234
rect 171 162 186 234
rect 284 162 299 234
<< ndiff >>
rect 36 96 65 106
rect 36 79 42 96
rect 59 79 65 96
rect 36 64 65 79
rect 80 96 109 106
rect 80 79 86 96
rect 103 79 109 96
rect 80 64 109 79
rect 142 96 171 106
rect 142 79 148 96
rect 165 79 171 96
rect 142 64 171 79
rect 186 96 215 106
rect 186 79 192 96
rect 209 79 215 96
rect 186 64 215 79
rect 255 96 284 106
rect 255 79 261 96
rect 278 79 284 96
rect 255 64 284 79
rect 299 96 328 106
rect 299 79 305 96
rect 322 79 328 96
rect 299 64 328 79
<< pdiff >>
rect 36 225 65 234
rect 36 208 42 225
rect 59 208 65 225
rect 36 191 65 208
rect 36 174 42 191
rect 59 174 65 191
rect 36 162 65 174
rect 80 217 109 234
rect 80 200 86 217
rect 103 200 109 217
rect 80 183 109 200
rect 80 166 86 183
rect 103 166 109 183
rect 80 162 109 166
rect 142 217 171 234
rect 142 200 148 217
rect 165 200 171 217
rect 142 183 171 200
rect 142 166 148 183
rect 165 166 171 183
rect 142 162 171 166
rect 186 217 215 234
rect 186 200 192 217
rect 209 200 215 217
rect 186 183 215 200
rect 186 166 192 183
rect 209 166 215 183
rect 186 162 215 166
rect 255 217 284 234
rect 255 200 261 217
rect 278 200 284 217
rect 255 183 284 200
rect 255 166 261 183
rect 278 166 284 183
rect 255 162 284 166
rect 299 217 328 234
rect 299 200 305 217
rect 322 200 328 217
rect 299 183 328 200
rect 299 166 305 183
rect 322 166 328 183
rect 299 162 328 166
<< ndiffc >>
rect 42 79 59 96
rect 86 79 103 96
rect 148 79 165 96
rect 192 79 209 96
rect 261 79 278 96
rect 305 79 322 96
<< pdiffc >>
rect 42 208 59 225
rect 42 174 59 191
rect 86 200 103 217
rect 86 166 103 183
rect 148 200 165 217
rect 148 166 165 183
rect 192 200 209 217
rect 192 166 209 183
rect 261 200 278 217
rect 261 166 278 183
rect 305 200 322 217
rect 305 166 322 183
<< psubdiff >>
rect 30 3 71 4
rect 30 -14 42 3
rect 59 -14 71 3
rect 30 -15 71 -14
<< nsubdiff >>
rect 30 279 72 280
rect 30 262 42 279
rect 59 262 72 279
rect 30 261 72 262
<< psubdiffcont >>
rect 42 -14 59 3
<< nsubdiffcont >>
rect 42 262 59 279
<< poly >>
rect 163 280 196 285
rect 163 263 171 280
rect 188 263 196 280
rect 163 258 196 263
rect 276 280 309 285
rect 276 263 284 280
rect 301 263 309 280
rect 276 258 309 263
rect 65 234 80 247
rect 171 234 186 258
rect 284 234 299 258
rect 65 106 80 162
rect 171 149 186 162
rect 284 149 299 162
rect 171 106 186 119
rect 284 106 299 119
rect 65 50 80 64
rect 171 50 186 64
rect 284 50 299 64
rect 65 45 110 50
rect 65 28 84 45
rect 101 28 110 45
rect 65 23 110 28
rect 163 45 196 50
rect 163 28 171 45
rect 188 28 196 45
rect 163 23 196 28
rect 276 45 309 50
rect 276 28 284 45
rect 301 28 309 45
rect 276 23 309 28
<< polycont >>
rect 171 263 188 280
rect 284 263 301 280
rect 84 28 101 45
rect 171 28 188 45
rect 284 28 301 45
<< locali >>
rect 42 279 59 293
rect 42 225 59 262
rect 42 191 59 208
rect 42 162 59 174
rect 86 280 244 282
rect 86 263 171 280
rect 188 263 244 280
rect 276 263 284 280
rect 301 263 309 280
rect 86 261 244 263
rect 86 217 103 261
rect 86 183 103 200
rect 42 96 59 106
rect 42 5 59 79
rect 86 96 103 166
rect 148 217 165 234
rect 148 183 165 200
rect 148 149 165 166
rect 133 143 165 149
rect 133 126 135 143
rect 152 126 165 143
rect 133 122 165 126
rect 86 70 103 79
rect 148 96 165 122
rect 148 70 165 79
rect 192 217 209 234
rect 192 183 209 200
rect 192 145 209 166
rect 192 96 209 128
rect 192 70 209 79
rect 227 48 244 261
rect 261 229 278 234
rect 261 183 278 200
rect 261 96 278 166
rect 261 70 278 79
rect 305 232 322 234
rect 305 229 334 232
rect 305 217 314 229
rect 331 212 334 229
rect 322 209 334 212
rect 305 183 322 200
rect 305 96 322 166
rect 305 70 322 79
rect 163 45 196 47
rect 76 28 84 45
rect 101 28 109 45
rect 163 28 171 45
rect 188 28 196 45
rect 163 26 196 28
rect 227 45 309 48
rect 227 28 284 45
rect 301 28 309 45
rect 227 27 309 28
rect 29 3 72 5
rect 29 -14 42 3
rect 59 -14 72 3
rect 29 -15 72 -14
<< viali >>
rect 284 263 301 280
rect 135 126 152 143
rect 192 128 209 145
rect 261 217 278 229
rect 261 212 278 217
rect 314 217 331 229
rect 314 212 322 217
rect 322 212 331 217
rect 84 28 101 45
rect 171 28 188 45
<< metal1 >>
rect 276 284 308 287
rect 276 258 279 284
rect 305 258 308 284
rect 276 255 308 258
rect 0 229 284 235
rect 0 212 261 229
rect 278 212 284 229
rect 0 206 284 212
rect 308 229 390 235
rect 308 212 314 229
rect 331 212 390 229
rect 308 206 390 212
rect 363 188 390 206
rect 363 151 408 188
rect 0 143 158 150
rect 0 126 135 143
rect 152 126 158 143
rect 0 120 158 126
rect 186 146 408 151
rect 186 145 392 146
rect 186 128 192 145
rect 209 128 392 145
rect 186 122 392 128
rect 163 51 195 52
rect 0 49 195 51
rect 0 45 166 49
rect 0 28 84 45
rect 101 28 166 45
rect 0 23 166 28
rect 192 23 195 49
rect 0 21 195 23
rect 163 20 195 21
<< via1 >>
rect 279 280 305 284
rect 279 263 284 280
rect 284 263 301 280
rect 301 263 305 280
rect 279 258 305 263
rect 166 45 192 49
rect 166 28 171 45
rect 171 28 188 45
rect 188 28 192 45
rect 166 23 192 28
<< metal2 >>
rect 276 284 308 287
rect 276 283 279 284
rect 223 258 279 283
rect 305 258 308 284
rect 163 51 195 52
rect 223 51 248 258
rect 276 255 308 258
rect 163 49 248 51
rect 163 23 166 49
rect 192 23 248 49
rect 163 21 248 23
rect 163 20 195 21
<< labels >>
rlabel metal1 s 0 36 0 36 4 SEL
port 1 nsew
rlabel metal1 s 0 220 0 220 4 A
port 2 nsew
rlabel metal1 s 0 135 0 135 4 B
port 3 nsew
rlabel metal1 s 408 167 408 167 4 Out
port 4 nsew
rlabel locali s 50 293 50 293 4 VDD
port 5 nsew
rlabel locali s 50 -3 50 -3 4 GND
port 6 nsew
<< end >>
