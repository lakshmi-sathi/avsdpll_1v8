magic
tech sky130A
magscale 1 2
timestamp 1607692587
<< nwell >>
rect -200 1928 30 1930
rect -200 1780 2980 1928
rect -200 96 3244 1780
rect -200 -56 2980 96
rect -200 -58 30 -56
<< nsubdiff >>
rect 110 1868 198 1872
rect 110 1834 134 1868
rect 168 1834 198 1868
rect 350 1868 438 1872
rect 350 1834 374 1868
rect 408 1834 438 1868
rect 590 1868 678 1872
rect 590 1834 614 1868
rect 648 1834 678 1868
rect 830 1868 918 1872
rect 830 1834 854 1868
rect 888 1834 918 1868
rect 1070 1868 1158 1872
rect 1070 1834 1094 1868
rect 1128 1834 1158 1868
rect 1310 1868 1398 1872
rect 1310 1834 1334 1868
rect 1368 1834 1398 1868
rect 1550 1868 1638 1872
rect 1550 1834 1574 1868
rect 1608 1834 1638 1868
rect 1790 1868 1878 1872
rect 1790 1834 1814 1868
rect 1848 1834 1878 1868
rect 2030 1868 2118 1872
rect 2030 1834 2054 1868
rect 2088 1834 2118 1868
rect 2270 1868 2358 1872
rect 2270 1834 2294 1868
rect 2328 1834 2358 1868
rect 2510 1868 2598 1872
rect 2510 1834 2534 1868
rect 2568 1834 2598 1868
rect 2750 1868 2838 1872
rect 2750 1834 2774 1868
rect 2808 1834 2838 1868
rect 108 42 196 46
rect 108 8 133 42
rect 167 8 196 42
rect 348 42 436 46
rect 348 8 373 42
rect 407 8 436 42
rect 588 42 676 46
rect 588 8 613 42
rect 647 8 676 42
rect 828 42 916 46
rect 828 8 853 42
rect 887 8 916 42
rect 1068 42 1156 46
rect 1068 8 1093 42
rect 1127 8 1156 42
rect 1308 42 1396 46
rect 1308 8 1333 42
rect 1367 8 1396 42
rect 1548 42 1636 46
rect 1548 8 1573 42
rect 1607 8 1636 42
rect 1788 42 1876 46
rect 1788 8 1813 42
rect 1847 8 1876 42
rect 2028 42 2116 46
rect 2028 8 2053 42
rect 2087 8 2116 42
rect 2268 42 2356 46
rect 2268 8 2293 42
rect 2327 8 2356 42
rect 2508 42 2596 46
rect 2508 8 2533 42
rect 2567 8 2596 42
rect 2748 42 2836 46
rect 2748 8 2773 42
rect 2807 8 2836 42
<< nsubdiffcont >>
rect 134 1834 168 1868
rect 374 1834 408 1868
rect 614 1834 648 1868
rect 854 1834 888 1868
rect 1094 1834 1128 1868
rect 1334 1834 1368 1868
rect 1574 1834 1608 1868
rect 1814 1834 1848 1868
rect 2054 1834 2088 1868
rect 2294 1834 2328 1868
rect 2534 1834 2568 1868
rect 2774 1834 2808 1868
rect 133 8 167 42
rect 373 8 407 42
rect 613 8 647 42
rect 853 8 887 42
rect 1093 8 1127 42
rect 1333 8 1367 42
rect 1573 8 1607 42
rect 1813 8 1847 42
rect 2053 8 2087 42
rect 2293 8 2327 42
rect 2533 8 2567 42
rect 2773 8 2807 42
<< locali >>
rect -24 1871 2956 1892
rect -24 1837 13 1871
rect 47 1868 253 1871
rect 47 1837 134 1868
rect -24 1834 134 1837
rect 168 1837 253 1868
rect 287 1868 493 1871
rect 287 1837 374 1868
rect 168 1834 374 1837
rect 408 1837 493 1868
rect 527 1868 733 1871
rect 527 1837 614 1868
rect 408 1834 614 1837
rect 648 1837 733 1868
rect 767 1868 973 1871
rect 767 1837 854 1868
rect 648 1834 854 1837
rect 888 1837 973 1868
rect 1007 1868 1213 1871
rect 1007 1837 1094 1868
rect 888 1834 1094 1837
rect 1128 1837 1213 1868
rect 1247 1868 1453 1871
rect 1247 1837 1334 1868
rect 1128 1834 1334 1837
rect 1368 1837 1453 1868
rect 1487 1868 1693 1871
rect 1487 1837 1574 1868
rect 1368 1834 1574 1837
rect 1608 1837 1693 1868
rect 1727 1868 1933 1871
rect 1727 1837 1814 1868
rect 1608 1834 1814 1837
rect 1848 1837 1933 1868
rect 1967 1868 2173 1871
rect 1967 1837 2054 1868
rect 1848 1834 2054 1837
rect 2088 1837 2173 1868
rect 2207 1868 2413 1871
rect 2207 1837 2294 1868
rect 2088 1834 2294 1837
rect 2328 1837 2413 1868
rect 2447 1868 2653 1871
rect 2447 1837 2534 1868
rect 2328 1834 2534 1837
rect 2568 1837 2653 1868
rect 2687 1868 2893 1871
rect 2687 1837 2774 1868
rect 2568 1834 2774 1837
rect 2808 1837 2893 1868
rect 2927 1837 2956 1871
rect 2808 1834 2956 1837
rect -24 1806 2956 1834
rect -130 986 -50 1348
rect -10 1026 70 1806
rect 110 986 190 1766
rect 230 1026 310 1806
rect 350 986 430 1766
rect 470 1026 550 1806
rect 590 986 670 1766
rect 710 1026 790 1806
rect 830 986 910 1766
rect 950 1026 1030 1806
rect 1070 986 1150 1766
rect 1190 1026 1270 1806
rect 1310 986 1390 1766
rect 1430 1026 1510 1806
rect 1550 986 1630 1766
rect 1670 1026 1750 1806
rect 1790 986 1870 1766
rect 1910 1026 1990 1806
rect 2030 986 2110 1766
rect 2150 1026 2230 1806
rect 2270 986 2350 1766
rect 2390 1026 2470 1806
rect 2510 986 2590 1766
rect 2630 1026 2710 1806
rect 2750 986 2830 1766
rect 2870 1026 2950 1806
rect 2990 986 3070 1766
rect 3134 986 3214 1368
rect -162 955 3244 986
rect -162 921 -107 955
rect -73 921 133 955
rect 167 921 373 955
rect 407 921 613 955
rect 647 921 853 955
rect 887 921 1093 955
rect 1127 921 1333 955
rect 1367 921 1573 955
rect 1607 921 1813 955
rect 1847 921 2053 955
rect 2087 921 2293 955
rect 2327 921 2533 955
rect 2567 921 2773 955
rect 2807 921 3013 955
rect 3047 921 3157 955
rect 3191 921 3244 955
rect -162 890 3244 921
rect -130 502 -50 890
rect -130 494 -60 502
rect -10 70 70 850
rect 110 110 190 890
rect 230 70 310 850
rect 350 110 430 890
rect 470 70 550 850
rect 590 110 670 890
rect 710 70 790 850
rect 830 110 910 890
rect 950 70 1030 850
rect 1070 110 1150 890
rect 1190 70 1270 850
rect 1310 110 1390 890
rect 1430 70 1510 850
rect 1550 110 1630 890
rect 1670 70 1750 850
rect 1790 110 1870 890
rect 1910 70 1990 850
rect 2030 110 2110 890
rect 2150 70 2230 850
rect 2270 110 2350 890
rect 2390 70 2470 850
rect 2510 110 2590 890
rect 2630 70 2710 850
rect 2750 110 2830 890
rect 2870 70 2950 850
rect 2990 110 3070 890
rect 3134 574 3214 890
rect -30 42 2956 70
rect -30 39 133 42
rect -30 5 13 39
rect 47 8 133 39
rect 167 39 373 42
rect 167 8 253 39
rect 47 5 253 8
rect 287 8 373 39
rect 407 39 613 42
rect 407 8 493 39
rect 287 5 493 8
rect 527 8 613 39
rect 647 39 853 42
rect 647 8 733 39
rect 527 5 733 8
rect 767 8 853 39
rect 887 39 1093 42
rect 887 8 973 39
rect 767 5 973 8
rect 1007 8 1093 39
rect 1127 39 1333 42
rect 1127 8 1213 39
rect 1007 5 1213 8
rect 1247 8 1333 39
rect 1367 39 1573 42
rect 1367 8 1453 39
rect 1247 5 1453 8
rect 1487 8 1573 39
rect 1607 39 1813 42
rect 1607 8 1693 39
rect 1487 5 1693 8
rect 1727 8 1813 39
rect 1847 39 2053 42
rect 1847 8 1933 39
rect 1727 5 1933 8
rect 1967 8 2053 39
rect 2087 39 2293 42
rect 2087 8 2173 39
rect 1967 5 2173 8
rect 2207 8 2293 39
rect 2327 39 2533 42
rect 2327 8 2413 39
rect 2207 5 2413 8
rect 2447 8 2533 39
rect 2567 39 2773 42
rect 2567 8 2653 39
rect 2447 5 2653 8
rect 2687 8 2773 39
rect 2807 39 2956 42
rect 2807 8 2893 39
rect 2687 5 2893 8
rect 2927 5 2956 39
rect -30 -16 2956 5
<< viali >>
rect 13 1837 47 1871
rect 253 1837 287 1871
rect 493 1837 527 1871
rect 733 1837 767 1871
rect 973 1837 1007 1871
rect 1213 1837 1247 1871
rect 1453 1837 1487 1871
rect 1693 1837 1727 1871
rect 1933 1837 1967 1871
rect 2173 1837 2207 1871
rect 2413 1837 2447 1871
rect 2653 1837 2687 1871
rect 2893 1837 2927 1871
rect -107 921 -73 955
rect 133 921 167 955
rect 373 921 407 955
rect 613 921 647 955
rect 853 921 887 955
rect 1093 921 1127 955
rect 1333 921 1367 955
rect 1573 921 1607 955
rect 1813 921 1847 955
rect 2053 921 2087 955
rect 2293 921 2327 955
rect 2533 921 2567 955
rect 2773 921 2807 955
rect 3013 921 3047 955
rect 3157 921 3191 955
rect 13 5 47 39
rect 253 5 287 39
rect 493 5 527 39
rect 733 5 767 39
rect 973 5 1007 39
rect 1213 5 1247 39
rect 1453 5 1487 39
rect 1693 5 1727 39
rect 1933 5 1967 39
rect 2173 5 2207 39
rect 2413 5 2447 39
rect 2653 5 2687 39
rect 2893 5 2927 39
<< metal1 >>
rect -24 1880 2956 1892
rect -24 1828 4 1880
rect 56 1828 244 1880
rect 296 1828 484 1880
rect 536 1828 724 1880
rect 776 1828 964 1880
rect 1016 1828 1204 1880
rect 1256 1828 1444 1880
rect 1496 1828 1684 1880
rect 1736 1828 1924 1880
rect 1976 1828 2164 1880
rect 2216 1828 2404 1880
rect 2456 1828 2644 1880
rect 2696 1828 2884 1880
rect 2936 1828 2956 1880
rect -24 1800 2956 1828
rect -136 992 -44 1348
rect -16 1020 76 1800
rect 104 992 196 1772
rect 224 1020 316 1800
rect 344 992 436 1772
rect 464 1020 556 1800
rect 584 992 676 1772
rect 704 1020 796 1800
rect 824 992 916 1772
rect 944 1020 1036 1800
rect 1064 992 1156 1772
rect 1184 1020 1276 1800
rect 1304 992 1396 1772
rect 1424 1020 1516 1800
rect 1544 992 1636 1772
rect 1664 1020 1756 1800
rect 1784 992 1876 1772
rect 1904 1020 1996 1800
rect 2024 992 2116 1772
rect 2144 1020 2236 1800
rect 2264 992 2356 1772
rect 2384 1020 2476 1800
rect 2504 992 2596 1772
rect 2624 1020 2716 1800
rect 2744 992 2836 1772
rect 2864 1020 2956 1800
rect 2984 992 3076 1772
rect 3128 992 3220 1368
rect -162 964 3244 992
rect -162 912 -116 964
rect -64 912 124 964
rect 176 912 364 964
rect 416 912 604 964
rect 656 912 844 964
rect 896 912 1084 964
rect 1136 912 1324 964
rect 1376 912 1564 964
rect 1616 912 1804 964
rect 1856 912 2044 964
rect 2096 912 2284 964
rect 2336 912 2524 964
rect 2576 912 2764 964
rect 2816 912 3004 964
rect 3056 912 3148 964
rect 3200 912 3244 964
rect -162 884 3244 912
rect -136 502 -44 884
rect -136 494 -60 502
rect -16 76 76 856
rect 104 104 196 884
rect 224 76 316 856
rect 344 104 436 884
rect 464 76 556 856
rect 584 104 676 884
rect 704 76 796 856
rect 824 104 916 884
rect 944 76 1036 856
rect 1064 104 1156 884
rect 1184 76 1276 856
rect 1304 104 1396 884
rect 1424 76 1516 856
rect 1544 104 1636 884
rect 1664 76 1756 856
rect 1784 104 1876 884
rect 1904 76 1996 856
rect 2024 104 2116 884
rect 2144 76 2236 856
rect 2264 104 2356 884
rect 2384 76 2476 856
rect 2504 104 2596 884
rect 2624 76 2716 856
rect 2744 104 2836 884
rect 2864 76 2956 856
rect 2984 104 3076 884
rect 3128 574 3220 884
rect -30 48 2956 76
rect -30 -4 4 48
rect 56 -4 244 48
rect 296 -4 484 48
rect 536 -4 724 48
rect 776 -4 964 48
rect 1016 -4 1204 48
rect 1256 -4 1444 48
rect 1496 -4 1684 48
rect 1736 -4 1924 48
rect 1976 -4 2164 48
rect 2216 -4 2404 48
rect 2456 -4 2644 48
rect 2696 -4 2884 48
rect 2936 -4 2956 48
rect -30 -16 2956 -4
<< via1 >>
rect 4 1871 56 1880
rect 4 1837 13 1871
rect 13 1837 47 1871
rect 47 1837 56 1871
rect 4 1828 56 1837
rect 244 1871 296 1880
rect 244 1837 253 1871
rect 253 1837 287 1871
rect 287 1837 296 1871
rect 244 1828 296 1837
rect 484 1871 536 1880
rect 484 1837 493 1871
rect 493 1837 527 1871
rect 527 1837 536 1871
rect 484 1828 536 1837
rect 724 1871 776 1880
rect 724 1837 733 1871
rect 733 1837 767 1871
rect 767 1837 776 1871
rect 724 1828 776 1837
rect 964 1871 1016 1880
rect 964 1837 973 1871
rect 973 1837 1007 1871
rect 1007 1837 1016 1871
rect 964 1828 1016 1837
rect 1204 1871 1256 1880
rect 1204 1837 1213 1871
rect 1213 1837 1247 1871
rect 1247 1837 1256 1871
rect 1204 1828 1256 1837
rect 1444 1871 1496 1880
rect 1444 1837 1453 1871
rect 1453 1837 1487 1871
rect 1487 1837 1496 1871
rect 1444 1828 1496 1837
rect 1684 1871 1736 1880
rect 1684 1837 1693 1871
rect 1693 1837 1727 1871
rect 1727 1837 1736 1871
rect 1684 1828 1736 1837
rect 1924 1871 1976 1880
rect 1924 1837 1933 1871
rect 1933 1837 1967 1871
rect 1967 1837 1976 1871
rect 1924 1828 1976 1837
rect 2164 1871 2216 1880
rect 2164 1837 2173 1871
rect 2173 1837 2207 1871
rect 2207 1837 2216 1871
rect 2164 1828 2216 1837
rect 2404 1871 2456 1880
rect 2404 1837 2413 1871
rect 2413 1837 2447 1871
rect 2447 1837 2456 1871
rect 2404 1828 2456 1837
rect 2644 1871 2696 1880
rect 2644 1837 2653 1871
rect 2653 1837 2687 1871
rect 2687 1837 2696 1871
rect 2644 1828 2696 1837
rect 2884 1871 2936 1880
rect 2884 1837 2893 1871
rect 2893 1837 2927 1871
rect 2927 1837 2936 1871
rect 2884 1828 2936 1837
rect -116 955 -64 964
rect -116 921 -107 955
rect -107 921 -73 955
rect -73 921 -64 955
rect -116 912 -64 921
rect 124 955 176 964
rect 124 921 133 955
rect 133 921 167 955
rect 167 921 176 955
rect 124 912 176 921
rect 364 955 416 964
rect 364 921 373 955
rect 373 921 407 955
rect 407 921 416 955
rect 364 912 416 921
rect 604 955 656 964
rect 604 921 613 955
rect 613 921 647 955
rect 647 921 656 955
rect 604 912 656 921
rect 844 955 896 964
rect 844 921 853 955
rect 853 921 887 955
rect 887 921 896 955
rect 844 912 896 921
rect 1084 955 1136 964
rect 1084 921 1093 955
rect 1093 921 1127 955
rect 1127 921 1136 955
rect 1084 912 1136 921
rect 1324 955 1376 964
rect 1324 921 1333 955
rect 1333 921 1367 955
rect 1367 921 1376 955
rect 1324 912 1376 921
rect 1564 955 1616 964
rect 1564 921 1573 955
rect 1573 921 1607 955
rect 1607 921 1616 955
rect 1564 912 1616 921
rect 1804 955 1856 964
rect 1804 921 1813 955
rect 1813 921 1847 955
rect 1847 921 1856 955
rect 1804 912 1856 921
rect 2044 955 2096 964
rect 2044 921 2053 955
rect 2053 921 2087 955
rect 2087 921 2096 955
rect 2044 912 2096 921
rect 2284 955 2336 964
rect 2284 921 2293 955
rect 2293 921 2327 955
rect 2327 921 2336 955
rect 2284 912 2336 921
rect 2524 955 2576 964
rect 2524 921 2533 955
rect 2533 921 2567 955
rect 2567 921 2576 955
rect 2524 912 2576 921
rect 2764 955 2816 964
rect 2764 921 2773 955
rect 2773 921 2807 955
rect 2807 921 2816 955
rect 2764 912 2816 921
rect 3004 955 3056 964
rect 3004 921 3013 955
rect 3013 921 3047 955
rect 3047 921 3056 955
rect 3004 912 3056 921
rect 3148 955 3200 964
rect 3148 921 3157 955
rect 3157 921 3191 955
rect 3191 921 3200 955
rect 3148 912 3200 921
rect 4 39 56 48
rect 4 5 13 39
rect 13 5 47 39
rect 47 5 56 39
rect 4 -4 56 5
rect 244 39 296 48
rect 244 5 253 39
rect 253 5 287 39
rect 287 5 296 39
rect 244 -4 296 5
rect 484 39 536 48
rect 484 5 493 39
rect 493 5 527 39
rect 527 5 536 39
rect 484 -4 536 5
rect 724 39 776 48
rect 724 5 733 39
rect 733 5 767 39
rect 767 5 776 39
rect 724 -4 776 5
rect 964 39 1016 48
rect 964 5 973 39
rect 973 5 1007 39
rect 1007 5 1016 39
rect 964 -4 1016 5
rect 1204 39 1256 48
rect 1204 5 1213 39
rect 1213 5 1247 39
rect 1247 5 1256 39
rect 1204 -4 1256 5
rect 1444 39 1496 48
rect 1444 5 1453 39
rect 1453 5 1487 39
rect 1487 5 1496 39
rect 1444 -4 1496 5
rect 1684 39 1736 48
rect 1684 5 1693 39
rect 1693 5 1727 39
rect 1727 5 1736 39
rect 1684 -4 1736 5
rect 1924 39 1976 48
rect 1924 5 1933 39
rect 1933 5 1967 39
rect 1967 5 1976 39
rect 1924 -4 1976 5
rect 2164 39 2216 48
rect 2164 5 2173 39
rect 2173 5 2207 39
rect 2207 5 2216 39
rect 2164 -4 2216 5
rect 2404 39 2456 48
rect 2404 5 2413 39
rect 2413 5 2447 39
rect 2447 5 2456 39
rect 2404 -4 2456 5
rect 2644 39 2696 48
rect 2644 5 2653 39
rect 2653 5 2687 39
rect 2687 5 2696 39
rect 2644 -4 2696 5
rect 2884 39 2936 48
rect 2884 5 2893 39
rect 2893 5 2927 39
rect 2927 5 2936 39
rect 2884 -4 2936 5
<< metal2 >>
rect -24 1882 2956 1892
rect -24 1826 2 1882
rect 58 1826 242 1882
rect 298 1826 482 1882
rect 538 1826 722 1882
rect 778 1826 962 1882
rect 1018 1826 1202 1882
rect 1258 1826 1442 1882
rect 1498 1826 1682 1882
rect 1738 1826 1922 1882
rect 1978 1826 2162 1882
rect 2218 1826 2402 1882
rect 2458 1826 2642 1882
rect 2698 1826 2882 1882
rect 2938 1826 2956 1882
rect -24 1800 2956 1826
rect -136 992 -44 1348
rect -16 1020 76 1800
rect 104 992 196 1772
rect 224 1020 316 1800
rect 344 992 436 1772
rect 464 1020 556 1800
rect 584 992 676 1772
rect 704 1020 796 1800
rect 824 992 916 1772
rect 944 1020 1036 1800
rect 1064 992 1156 1772
rect 1184 1020 1276 1800
rect 1304 992 1396 1772
rect 1424 1020 1516 1800
rect 1544 992 1636 1772
rect 1664 1020 1756 1800
rect 1784 992 1876 1772
rect 1904 1020 1996 1800
rect 2024 992 2116 1772
rect 2144 1020 2236 1800
rect 2264 992 2356 1772
rect 2384 1020 2476 1800
rect 2504 992 2596 1772
rect 2624 1020 2716 1800
rect 2744 992 2836 1772
rect 2864 1020 2956 1800
rect 2984 992 3076 1772
rect 3128 992 3220 1368
rect -162 966 3244 992
rect -162 910 -118 966
rect -62 910 122 966
rect 178 910 362 966
rect 418 910 602 966
rect 658 910 842 966
rect 898 910 1082 966
rect 1138 910 1322 966
rect 1378 910 1562 966
rect 1618 910 1802 966
rect 1858 910 2042 966
rect 2098 910 2282 966
rect 2338 910 2522 966
rect 2578 910 2762 966
rect 2818 910 3002 966
rect 3058 910 3146 966
rect 3202 910 3244 966
rect -162 884 3244 910
rect -136 502 -44 884
rect -136 494 -60 502
rect -16 76 76 856
rect 104 104 196 884
rect 224 76 316 856
rect 344 104 436 884
rect 464 76 556 856
rect 584 104 676 884
rect 704 76 796 856
rect 824 104 916 884
rect 944 76 1036 856
rect 1064 104 1156 884
rect 1184 76 1276 856
rect 1304 104 1396 884
rect 1424 76 1516 856
rect 1544 104 1636 884
rect 1664 76 1756 856
rect 1784 104 1876 884
rect 1904 76 1996 856
rect 2024 104 2116 884
rect 2144 76 2236 856
rect 2264 104 2356 884
rect 2384 76 2476 856
rect 2504 104 2596 884
rect 2624 76 2716 856
rect 2744 104 2836 884
rect 2864 76 2956 856
rect 2984 104 3076 884
rect 3128 574 3220 884
rect -30 50 2956 76
rect -30 -6 2 50
rect 58 -6 242 50
rect 298 -6 482 50
rect 538 -6 722 50
rect 778 -6 962 50
rect 1018 -6 1202 50
rect 1258 -6 1442 50
rect 1498 -6 1682 50
rect 1738 -6 1922 50
rect 1978 -6 2162 50
rect 2218 -6 2402 50
rect 2458 -6 2642 50
rect 2698 -6 2882 50
rect 2938 -6 2956 50
rect -30 -16 2956 -6
<< via2 >>
rect 2 1880 58 1882
rect 2 1828 4 1880
rect 4 1828 56 1880
rect 56 1828 58 1880
rect 2 1826 58 1828
rect 242 1880 298 1882
rect 242 1828 244 1880
rect 244 1828 296 1880
rect 296 1828 298 1880
rect 242 1826 298 1828
rect 482 1880 538 1882
rect 482 1828 484 1880
rect 484 1828 536 1880
rect 536 1828 538 1880
rect 482 1826 538 1828
rect 722 1880 778 1882
rect 722 1828 724 1880
rect 724 1828 776 1880
rect 776 1828 778 1880
rect 722 1826 778 1828
rect 962 1880 1018 1882
rect 962 1828 964 1880
rect 964 1828 1016 1880
rect 1016 1828 1018 1880
rect 962 1826 1018 1828
rect 1202 1880 1258 1882
rect 1202 1828 1204 1880
rect 1204 1828 1256 1880
rect 1256 1828 1258 1880
rect 1202 1826 1258 1828
rect 1442 1880 1498 1882
rect 1442 1828 1444 1880
rect 1444 1828 1496 1880
rect 1496 1828 1498 1880
rect 1442 1826 1498 1828
rect 1682 1880 1738 1882
rect 1682 1828 1684 1880
rect 1684 1828 1736 1880
rect 1736 1828 1738 1880
rect 1682 1826 1738 1828
rect 1922 1880 1978 1882
rect 1922 1828 1924 1880
rect 1924 1828 1976 1880
rect 1976 1828 1978 1880
rect 1922 1826 1978 1828
rect 2162 1880 2218 1882
rect 2162 1828 2164 1880
rect 2164 1828 2216 1880
rect 2216 1828 2218 1880
rect 2162 1826 2218 1828
rect 2402 1880 2458 1882
rect 2402 1828 2404 1880
rect 2404 1828 2456 1880
rect 2456 1828 2458 1880
rect 2402 1826 2458 1828
rect 2642 1880 2698 1882
rect 2642 1828 2644 1880
rect 2644 1828 2696 1880
rect 2696 1828 2698 1880
rect 2642 1826 2698 1828
rect 2882 1880 2938 1882
rect 2882 1828 2884 1880
rect 2884 1828 2936 1880
rect 2936 1828 2938 1880
rect 2882 1826 2938 1828
rect -118 964 -62 966
rect -118 912 -116 964
rect -116 912 -64 964
rect -64 912 -62 964
rect -118 910 -62 912
rect 122 964 178 966
rect 122 912 124 964
rect 124 912 176 964
rect 176 912 178 964
rect 122 910 178 912
rect 362 964 418 966
rect 362 912 364 964
rect 364 912 416 964
rect 416 912 418 964
rect 362 910 418 912
rect 602 964 658 966
rect 602 912 604 964
rect 604 912 656 964
rect 656 912 658 964
rect 602 910 658 912
rect 842 964 898 966
rect 842 912 844 964
rect 844 912 896 964
rect 896 912 898 964
rect 842 910 898 912
rect 1082 964 1138 966
rect 1082 912 1084 964
rect 1084 912 1136 964
rect 1136 912 1138 964
rect 1082 910 1138 912
rect 1322 964 1378 966
rect 1322 912 1324 964
rect 1324 912 1376 964
rect 1376 912 1378 964
rect 1322 910 1378 912
rect 1562 964 1618 966
rect 1562 912 1564 964
rect 1564 912 1616 964
rect 1616 912 1618 964
rect 1562 910 1618 912
rect 1802 964 1858 966
rect 1802 912 1804 964
rect 1804 912 1856 964
rect 1856 912 1858 964
rect 1802 910 1858 912
rect 2042 964 2098 966
rect 2042 912 2044 964
rect 2044 912 2096 964
rect 2096 912 2098 964
rect 2042 910 2098 912
rect 2282 964 2338 966
rect 2282 912 2284 964
rect 2284 912 2336 964
rect 2336 912 2338 964
rect 2282 910 2338 912
rect 2522 964 2578 966
rect 2522 912 2524 964
rect 2524 912 2576 964
rect 2576 912 2578 964
rect 2522 910 2578 912
rect 2762 964 2818 966
rect 2762 912 2764 964
rect 2764 912 2816 964
rect 2816 912 2818 964
rect 2762 910 2818 912
rect 3002 964 3058 966
rect 3002 912 3004 964
rect 3004 912 3056 964
rect 3056 912 3058 964
rect 3002 910 3058 912
rect 3146 964 3202 966
rect 3146 912 3148 964
rect 3148 912 3200 964
rect 3200 912 3202 964
rect 3146 910 3202 912
rect 2 48 58 50
rect 2 -4 4 48
rect 4 -4 56 48
rect 56 -4 58 48
rect 2 -6 58 -4
rect 242 48 298 50
rect 242 -4 244 48
rect 244 -4 296 48
rect 296 -4 298 48
rect 242 -6 298 -4
rect 482 48 538 50
rect 482 -4 484 48
rect 484 -4 536 48
rect 536 -4 538 48
rect 482 -6 538 -4
rect 722 48 778 50
rect 722 -4 724 48
rect 724 -4 776 48
rect 776 -4 778 48
rect 722 -6 778 -4
rect 962 48 1018 50
rect 962 -4 964 48
rect 964 -4 1016 48
rect 1016 -4 1018 48
rect 962 -6 1018 -4
rect 1202 48 1258 50
rect 1202 -4 1204 48
rect 1204 -4 1256 48
rect 1256 -4 1258 48
rect 1202 -6 1258 -4
rect 1442 48 1498 50
rect 1442 -4 1444 48
rect 1444 -4 1496 48
rect 1496 -4 1498 48
rect 1442 -6 1498 -4
rect 1682 48 1738 50
rect 1682 -4 1684 48
rect 1684 -4 1736 48
rect 1736 -4 1738 48
rect 1682 -6 1738 -4
rect 1922 48 1978 50
rect 1922 -4 1924 48
rect 1924 -4 1976 48
rect 1976 -4 1978 48
rect 1922 -6 1978 -4
rect 2162 48 2218 50
rect 2162 -4 2164 48
rect 2164 -4 2216 48
rect 2216 -4 2218 48
rect 2162 -6 2218 -4
rect 2402 48 2458 50
rect 2402 -4 2404 48
rect 2404 -4 2456 48
rect 2456 -4 2458 48
rect 2402 -6 2458 -4
rect 2642 48 2698 50
rect 2642 -4 2644 48
rect 2644 -4 2696 48
rect 2696 -4 2698 48
rect 2642 -6 2698 -4
rect 2882 48 2938 50
rect 2882 -4 2884 48
rect 2884 -4 2936 48
rect 2936 -4 2938 48
rect 2882 -6 2938 -4
<< metal3 >>
rect -24 1886 2956 1892
rect -24 1822 -2 1886
rect 62 1822 238 1886
rect 302 1822 478 1886
rect 542 1822 718 1886
rect 782 1822 958 1886
rect 1022 1822 1198 1886
rect 1262 1822 1438 1886
rect 1502 1822 1678 1886
rect 1742 1822 1918 1886
rect 1982 1822 2158 1886
rect 2222 1822 2398 1886
rect 2462 1822 2638 1886
rect 2702 1822 2878 1886
rect 2942 1822 2956 1886
rect -24 1816 2956 1822
rect -120 976 -60 1348
rect 0 1036 60 1816
rect 120 976 180 1756
rect 240 1036 300 1816
rect 360 976 420 1756
rect 480 1036 540 1816
rect 600 976 660 1756
rect 720 1036 780 1816
rect 840 976 900 1756
rect 960 1036 1020 1816
rect 1080 976 1140 1756
rect 1200 1036 1260 1816
rect 1320 976 1380 1756
rect 1440 1036 1500 1816
rect 1560 976 1620 1756
rect 1680 1036 1740 1816
rect 1800 976 1860 1756
rect 1920 1036 1980 1816
rect 2040 976 2100 1756
rect 2160 1036 2220 1816
rect 2280 976 2340 1756
rect 2400 1036 2460 1816
rect 2520 976 2580 1756
rect 2640 1036 2700 1816
rect 2760 976 2820 1756
rect 2880 1036 2940 1816
rect 3000 976 3060 1756
rect 3144 976 3204 1368
rect -162 970 3244 976
rect -162 906 -122 970
rect -58 906 118 970
rect 182 906 358 970
rect 422 906 598 970
rect 662 906 838 970
rect 902 906 1078 970
rect 1142 906 1318 970
rect 1382 906 1558 970
rect 1622 906 1798 970
rect 1862 906 2038 970
rect 2102 906 2278 970
rect 2342 906 2518 970
rect 2582 906 2758 970
rect 2822 906 2998 970
rect 3062 906 3142 970
rect 3206 906 3244 970
rect -162 900 3244 906
rect -120 494 -60 900
rect 0 60 60 840
rect 120 120 180 900
rect 240 60 300 840
rect 360 120 420 900
rect 480 60 540 840
rect 600 120 660 900
rect 720 60 780 840
rect 840 120 900 900
rect 960 60 1020 840
rect 1080 120 1140 900
rect 1200 60 1260 840
rect 1320 120 1380 900
rect 1440 60 1500 840
rect 1560 120 1620 900
rect 1680 60 1740 840
rect 1800 120 1860 900
rect 1920 60 1980 840
rect 2040 120 2100 900
rect 2160 60 2220 840
rect 2280 120 2340 900
rect 2400 60 2460 840
rect 2520 120 2580 900
rect 2640 60 2700 840
rect 2760 120 2820 900
rect 2880 60 2940 840
rect 3000 120 3060 900
rect 3144 574 3204 900
rect -30 54 2956 60
rect -30 -10 -2 54
rect 62 -10 238 54
rect 302 -10 478 54
rect 542 -10 718 54
rect 782 -10 958 54
rect 1022 -10 1198 54
rect 1262 -10 1438 54
rect 1502 -10 1678 54
rect 1742 -10 1918 54
rect 1982 -10 2158 54
rect 2222 -10 2398 54
rect 2462 -10 2638 54
rect 2702 -10 2878 54
rect 2942 -10 2956 54
rect -30 -16 2956 -10
<< via3 >>
rect -2 1882 62 1886
rect -2 1826 2 1882
rect 2 1826 58 1882
rect 58 1826 62 1882
rect -2 1822 62 1826
rect 238 1882 302 1886
rect 238 1826 242 1882
rect 242 1826 298 1882
rect 298 1826 302 1882
rect 238 1822 302 1826
rect 478 1882 542 1886
rect 478 1826 482 1882
rect 482 1826 538 1882
rect 538 1826 542 1882
rect 478 1822 542 1826
rect 718 1882 782 1886
rect 718 1826 722 1882
rect 722 1826 778 1882
rect 778 1826 782 1882
rect 718 1822 782 1826
rect 958 1882 1022 1886
rect 958 1826 962 1882
rect 962 1826 1018 1882
rect 1018 1826 1022 1882
rect 958 1822 1022 1826
rect 1198 1882 1262 1886
rect 1198 1826 1202 1882
rect 1202 1826 1258 1882
rect 1258 1826 1262 1882
rect 1198 1822 1262 1826
rect 1438 1882 1502 1886
rect 1438 1826 1442 1882
rect 1442 1826 1498 1882
rect 1498 1826 1502 1882
rect 1438 1822 1502 1826
rect 1678 1882 1742 1886
rect 1678 1826 1682 1882
rect 1682 1826 1738 1882
rect 1738 1826 1742 1882
rect 1678 1822 1742 1826
rect 1918 1882 1982 1886
rect 1918 1826 1922 1882
rect 1922 1826 1978 1882
rect 1978 1826 1982 1882
rect 1918 1822 1982 1826
rect 2158 1882 2222 1886
rect 2158 1826 2162 1882
rect 2162 1826 2218 1882
rect 2218 1826 2222 1882
rect 2158 1822 2222 1826
rect 2398 1882 2462 1886
rect 2398 1826 2402 1882
rect 2402 1826 2458 1882
rect 2458 1826 2462 1882
rect 2398 1822 2462 1826
rect 2638 1882 2702 1886
rect 2638 1826 2642 1882
rect 2642 1826 2698 1882
rect 2698 1826 2702 1882
rect 2638 1822 2702 1826
rect 2878 1882 2942 1886
rect 2878 1826 2882 1882
rect 2882 1826 2938 1882
rect 2938 1826 2942 1882
rect 2878 1822 2942 1826
rect -122 966 -58 970
rect -122 910 -118 966
rect -118 910 -62 966
rect -62 910 -58 966
rect -122 906 -58 910
rect 118 966 182 970
rect 118 910 122 966
rect 122 910 178 966
rect 178 910 182 966
rect 118 906 182 910
rect 358 966 422 970
rect 358 910 362 966
rect 362 910 418 966
rect 418 910 422 966
rect 358 906 422 910
rect 598 966 662 970
rect 598 910 602 966
rect 602 910 658 966
rect 658 910 662 966
rect 598 906 662 910
rect 838 966 902 970
rect 838 910 842 966
rect 842 910 898 966
rect 898 910 902 966
rect 838 906 902 910
rect 1078 966 1142 970
rect 1078 910 1082 966
rect 1082 910 1138 966
rect 1138 910 1142 966
rect 1078 906 1142 910
rect 1318 966 1382 970
rect 1318 910 1322 966
rect 1322 910 1378 966
rect 1378 910 1382 966
rect 1318 906 1382 910
rect 1558 966 1622 970
rect 1558 910 1562 966
rect 1562 910 1618 966
rect 1618 910 1622 966
rect 1558 906 1622 910
rect 1798 966 1862 970
rect 1798 910 1802 966
rect 1802 910 1858 966
rect 1858 910 1862 966
rect 1798 906 1862 910
rect 2038 966 2102 970
rect 2038 910 2042 966
rect 2042 910 2098 966
rect 2098 910 2102 966
rect 2038 906 2102 910
rect 2278 966 2342 970
rect 2278 910 2282 966
rect 2282 910 2338 966
rect 2338 910 2342 966
rect 2278 906 2342 910
rect 2518 966 2582 970
rect 2518 910 2522 966
rect 2522 910 2578 966
rect 2578 910 2582 966
rect 2518 906 2582 910
rect 2758 966 2822 970
rect 2758 910 2762 966
rect 2762 910 2818 966
rect 2818 910 2822 966
rect 2758 906 2822 910
rect 2998 966 3062 970
rect 2998 910 3002 966
rect 3002 910 3058 966
rect 3058 910 3062 966
rect 2998 906 3062 910
rect 3142 966 3206 970
rect 3142 910 3146 966
rect 3146 910 3202 966
rect 3202 910 3206 966
rect 3142 906 3206 910
rect -2 50 62 54
rect -2 -6 2 50
rect 2 -6 58 50
rect 58 -6 62 50
rect -2 -10 62 -6
rect 238 50 302 54
rect 238 -6 242 50
rect 242 -6 298 50
rect 298 -6 302 50
rect 238 -10 302 -6
rect 478 50 542 54
rect 478 -6 482 50
rect 482 -6 538 50
rect 538 -6 542 50
rect 478 -10 542 -6
rect 718 50 782 54
rect 718 -6 722 50
rect 722 -6 778 50
rect 778 -6 782 50
rect 718 -10 782 -6
rect 958 50 1022 54
rect 958 -6 962 50
rect 962 -6 1018 50
rect 1018 -6 1022 50
rect 958 -10 1022 -6
rect 1198 50 1262 54
rect 1198 -6 1202 50
rect 1202 -6 1258 50
rect 1258 -6 1262 50
rect 1198 -10 1262 -6
rect 1438 50 1502 54
rect 1438 -6 1442 50
rect 1442 -6 1498 50
rect 1498 -6 1502 50
rect 1438 -10 1502 -6
rect 1678 50 1742 54
rect 1678 -6 1682 50
rect 1682 -6 1738 50
rect 1738 -6 1742 50
rect 1678 -10 1742 -6
rect 1918 50 1982 54
rect 1918 -6 1922 50
rect 1922 -6 1978 50
rect 1978 -6 1982 50
rect 1918 -10 1982 -6
rect 2158 50 2222 54
rect 2158 -6 2162 50
rect 2162 -6 2218 50
rect 2218 -6 2222 50
rect 2158 -10 2222 -6
rect 2398 50 2462 54
rect 2398 -6 2402 50
rect 2402 -6 2458 50
rect 2458 -6 2462 50
rect 2398 -10 2462 -6
rect 2638 50 2702 54
rect 2638 -6 2642 50
rect 2642 -6 2698 50
rect 2698 -6 2702 50
rect 2638 -10 2702 -6
rect 2878 50 2942 54
rect 2878 -6 2882 50
rect 2882 -6 2938 50
rect 2938 -6 2942 50
rect 2878 -10 2942 -6
<< metal4 >>
rect -24 1886 2956 1892
rect -24 1822 -2 1886
rect 62 1822 238 1886
rect 302 1822 478 1886
rect 542 1822 718 1886
rect 782 1822 958 1886
rect 1022 1822 1198 1886
rect 1262 1822 1438 1886
rect 1502 1822 1678 1886
rect 1742 1822 1918 1886
rect 1982 1822 2158 1886
rect 2222 1822 2398 1886
rect 2462 1822 2638 1886
rect 2702 1822 2878 1886
rect 2942 1822 2956 1886
rect -24 1816 2956 1822
rect -120 976 -60 1348
rect 0 1036 60 1816
rect 120 976 180 1756
rect 240 1036 300 1816
rect 360 976 420 1756
rect 480 1036 540 1816
rect 600 976 660 1756
rect 720 1036 780 1816
rect 840 976 900 1756
rect 960 1036 1020 1816
rect 1080 976 1140 1756
rect 1200 1036 1260 1816
rect 1320 976 1380 1756
rect 1440 1036 1500 1816
rect 1560 976 1620 1756
rect 1680 1036 1740 1816
rect 1800 976 1860 1756
rect 1920 1036 1980 1816
rect 2040 976 2100 1756
rect 2160 1036 2220 1816
rect 2280 976 2340 1756
rect 2400 1036 2460 1816
rect 2520 976 2580 1756
rect 2640 1036 2700 1816
rect 2760 976 2820 1756
rect 2880 1036 2940 1816
rect 3000 976 3060 1756
rect 3144 976 3204 1368
rect -162 970 3244 976
rect -162 906 -122 970
rect -58 906 118 970
rect 182 906 358 970
rect 422 906 598 970
rect 662 906 838 970
rect 902 906 1078 970
rect 1142 906 1318 970
rect 1382 906 1558 970
rect 1622 906 1798 970
rect 1862 906 2038 970
rect 2102 906 2278 970
rect 2342 906 2518 970
rect 2582 906 2758 970
rect 2822 906 2998 970
rect 3062 906 3142 970
rect 3206 906 3244 970
rect -162 900 3244 906
rect -120 494 -60 900
rect 0 60 60 840
rect 120 120 180 900
rect 240 60 300 840
rect 360 120 420 900
rect 480 60 540 840
rect 600 120 660 900
rect 720 60 780 840
rect 840 120 900 900
rect 960 60 1020 840
rect 1080 120 1140 900
rect 1200 60 1260 840
rect 1320 120 1380 900
rect 1440 60 1500 840
rect 1560 120 1620 900
rect 1680 60 1740 840
rect 1800 120 1860 900
rect 1920 60 1980 840
rect 2040 120 2100 900
rect 2160 60 2220 840
rect 2280 120 2340 900
rect 2400 60 2460 840
rect 2520 120 2580 900
rect 2640 60 2700 840
rect 2760 120 2820 900
rect 2880 60 2940 840
rect 3000 120 3060 900
rect 3144 574 3204 900
rect -30 54 2956 60
rect -30 -10 -2 54
rect 62 -10 238 54
rect 302 -10 478 54
rect 542 -10 718 54
rect 782 -10 958 54
rect 1022 -10 1198 54
rect 1262 -10 1438 54
rect 1502 -10 1678 54
rect 1742 -10 1918 54
rect 1982 -10 2158 54
rect 2222 -10 2398 54
rect 2462 -10 2638 54
rect 2702 -10 2878 54
rect 2942 -10 2956 54
rect -30 -16 2956 -10
<< labels >>
rlabel metal4 s 150 -16 150 -16 4 pin1
port 1 nsew
rlabel metal4 s 390 -16 390 -16 4 pin1
port 1 nsew
rlabel metal4 s 630 -16 630 -16 4 pin1
port 1 nsew
rlabel metal4 s 630 1892 630 1892 4 pin1
port 1 nsew
rlabel metal4 s 390 1892 390 1892 4 pin1
port 1 nsew
rlabel metal4 s 150 1892 150 1892 4 pin1
port 1 nsew
rlabel metal4 s 870 -16 870 -16 4 pin1
port 1 nsew
rlabel metal4 s 1110 -16 1110 -16 4 pin1
port 1 nsew
rlabel metal4 s 1350 -16 1350 -16 4 pin1
port 1 nsew
rlabel metal4 s 1350 1892 1350 1892 4 pin1
port 1 nsew
rlabel metal4 s 1110 1892 1110 1892 4 pin1
port 1 nsew
rlabel metal4 s 870 1892 870 1892 4 pin1
port 1 nsew
rlabel metal4 s 1590 -16 1590 -16 4 pin1
port 1 nsew
rlabel metal4 s 1830 -16 1830 -16 4 pin1
port 1 nsew
rlabel metal4 s 2070 -16 2070 -16 4 pin1
port 1 nsew
rlabel metal4 s 2070 1892 2070 1892 4 pin1
port 1 nsew
rlabel metal4 s 1830 1892 1830 1892 4 pin1
port 1 nsew
rlabel metal4 s 1590 1892 1590 1892 4 pin1
port 1 nsew
rlabel metal4 s 2310 -16 2310 -16 4 pin1
port 1 nsew
rlabel metal4 s 2550 -16 2550 -16 4 pin1
port 1 nsew
rlabel metal4 s 2790 -16 2790 -16 4 pin1
port 1 nsew
rlabel metal4 s 2790 1892 2790 1892 4 pin1
port 1 nsew
rlabel metal4 s 2550 1892 2550 1892 4 pin1
port 1 nsew
rlabel metal4 s 2310 1892 2310 1892 4 pin1
port 1 nsew
rlabel metal4 s 148 976 148 976 4 pin2
port 2 nsew
rlabel metal4 s 388 976 388 976 4 pin2
port 2 nsew
rlabel metal4 s 628 976 628 976 4 pin2
port 2 nsew
rlabel metal4 s 628 900 628 900 4 pin2
port 2 nsew
rlabel metal4 s 388 900 388 900 4 pin2
port 2 nsew
rlabel metal4 s 148 900 148 900 4 pin2
port 2 nsew
rlabel metal4 s 868 976 868 976 4 pin2
port 2 nsew
rlabel metal4 s 1108 976 1108 976 4 pin2
port 2 nsew
rlabel metal4 s 1348 976 1348 976 4 pin2
port 2 nsew
rlabel metal4 s 1348 900 1348 900 4 pin2
port 2 nsew
rlabel metal4 s 1108 900 1108 900 4 pin2
port 2 nsew
rlabel metal4 s 868 900 868 900 4 pin2
port 2 nsew
rlabel metal4 s 1588 976 1588 976 4 pin2
port 2 nsew
rlabel metal4 s 1828 976 1828 976 4 pin2
port 2 nsew
rlabel metal4 s 2068 976 2068 976 4 pin2
port 2 nsew
rlabel metal4 s 2068 900 2068 900 4 pin2
port 2 nsew
rlabel metal4 s 1828 900 1828 900 4 pin2
port 2 nsew
rlabel metal4 s 1588 900 1588 900 4 pin2
port 2 nsew
rlabel metal4 s 2308 976 2308 976 4 pin2
port 2 nsew
rlabel metal4 s 2548 976 2548 976 4 pin2
port 2 nsew
rlabel metal4 s 2788 976 2788 976 4 pin2
port 2 nsew
rlabel metal4 s 2788 900 2788 900 4 pin2
port 2 nsew
rlabel metal4 s 2548 900 2548 900 4 pin2
port 2 nsew
rlabel metal4 s 2308 900 2308 900 4 pin2
port 2 nsew
rlabel metal4 s 3028 976 3028 976 4 pin2
port 2 nsew
rlabel metal4 s 3028 900 3028 900 4 pin2
port 2 nsew
rlabel metal4 s 3172 900 3172 900 4 pin2
port 2 nsew
rlabel metal4 s 3172 976 3172 976 4 pin2
port 2 nsew
rlabel metal4 s -92 976 -92 976 4 pin2
port 2 nsew
rlabel metal4 s -92 900 -92 900 4 pin2
port 2 nsew
<< end >>
