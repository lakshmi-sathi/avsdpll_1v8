magic
tech sky130A
magscale 1 2
timestamp 1607692587
<< pwell >>
rect -175 215 175 249
rect -175 -215 -141 215
rect 141 -215 175 215
rect -175 -249 175 -215
<< nmos >>
rect -15 -75 15 75
<< ndiff >>
rect -73 51 -15 75
rect -73 17 -61 51
rect -27 17 -15 51
rect -73 -17 -15 17
rect -73 -51 -61 -17
rect -27 -51 -15 -17
rect -73 -75 -15 -51
rect 15 51 73 75
rect 15 17 27 51
rect 61 17 73 51
rect 15 -17 73 17
rect 15 -51 27 -17
rect 61 -51 73 -17
rect 15 -75 73 -51
<< ndiffc >>
rect -61 17 -27 51
rect -61 -51 -27 -17
rect 27 17 61 51
rect 27 -51 61 -17
<< psubdiff >>
rect -175 215 -51 249
rect -17 215 17 249
rect 51 215 175 249
rect -175 153 -141 215
rect -175 85 -141 119
rect 141 153 175 215
rect 141 85 175 119
rect -175 17 -141 51
rect -175 -51 -141 -17
rect 141 17 175 51
rect 141 -51 175 -17
rect -175 -119 -141 -85
rect -175 -215 -141 -153
rect 141 -119 175 -85
rect 141 -215 175 -153
rect -175 -249 -51 -215
rect -17 -249 17 -215
rect 51 -249 175 -215
<< psubdiffcont >>
rect -51 215 -17 249
rect 17 215 51 249
rect -175 119 -141 153
rect 141 119 175 153
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect -175 -153 -141 -119
rect 141 -153 175 -119
rect -51 -249 -17 -215
rect 17 -249 51 -215
<< poly >>
rect -69 151 69 167
rect -69 117 -53 151
rect -19 117 19 151
rect 53 117 69 151
rect -69 97 69 117
rect -15 75 15 97
rect -15 -97 15 -75
rect -33 -163 33 -97
<< polycont >>
rect -53 117 -19 151
rect 19 117 53 151
<< locali >>
rect -175 215 -51 249
rect -17 215 17 249
rect 51 215 175 249
rect -175 153 -141 215
rect 141 153 175 215
rect -175 85 -141 119
rect -69 117 -53 151
rect -19 117 19 151
rect 53 117 69 151
rect 141 85 175 119
rect -175 17 -141 51
rect -175 -51 -141 -17
rect -61 53 -27 79
rect -61 -17 -27 17
rect -61 -79 -27 -53
rect 27 53 61 79
rect 27 -17 61 17
rect 27 -79 61 -53
rect 141 17 175 51
rect 141 -51 175 -17
rect -175 -119 -141 -85
rect -175 -215 -141 -153
rect 141 -119 175 -85
rect 141 -215 175 -153
rect -175 -249 -51 -215
rect -17 -249 17 -215
rect 51 -249 175 -215
<< viali >>
rect -53 117 -19 151
rect 19 117 53 151
rect -61 51 -27 53
rect -61 19 -27 51
rect -61 -51 -27 -19
rect -61 -53 -27 -51
rect 27 51 61 53
rect 27 19 61 51
rect 27 -51 61 -19
rect 27 -53 61 -51
<< metal1 >>
rect -81 117 -71 169
rect -19 117 19 169
rect 71 117 81 169
rect -81 111 81 117
rect -67 53 -21 75
rect -67 19 -61 53
rect -27 19 -21 53
rect -67 -19 -21 19
rect -67 -53 -61 -19
rect -27 -53 -21 -19
rect -67 -75 -21 -53
rect 21 53 67 75
rect 21 19 27 53
rect 61 19 67 53
rect 21 -19 67 19
rect 21 -53 27 -19
rect 61 -53 67 -19
rect 21 -75 67 -53
<< via1 >>
rect -71 151 -19 169
rect -71 117 -53 151
rect -53 117 -19 151
rect 19 151 71 169
rect 19 117 53 151
rect 53 117 71 151
<< metal2 >>
rect -71 169 71 179
rect -19 117 19 169
rect -71 107 71 117
<< properties >>
string FIXED_BBOX -158 -232 158 232
<< end >>
