* SPICE3 file created from VCO_fin.ext - technology: sky130A
.include sky130nm.lib
.option scale=0.01u

XM1000 VDD a_n90_303# a_0_94# VDD sky130_fd_pr__pfet_01v8 w=108 l=15
+  ad=3132 pd=278.64 as=3132 ps=299.52
XM1001 a_144_n15# a_44_n15# a_0_94# VDD sky130_fd_pr__pfet_01v8 w=42 l=15
+  ad=1218 pd=142 as=1218 ps=116.48
XM1002 a_0_46# a_544_n15# a_0_n15# GND sky130_fd_pr__nfet_01v8 w=120 l=15
+  ad=3480 pd=298 as=3480 ps=356
XM1003 GND VCtrl a_0_n15# GND sky130_fd_pr__nfet_01v8 w=108 l=15
+  ad=3132 pd=292.39 as=3132 ps=320.4
XM1004 a_44_n15# a_0_46# a_0_94# VDD sky130_fd_pr__pfet_01v8 w=42 l=15
+  ad=1218 pd=142 as=1218 ps=116.48
XM1005 Clk_Out a_0_46# GND GND sky130_fd_pr__nfet_01v8 w=54 l=15
+  ad=1566 pd=166 as=1566 ps=146.195
XM1006 a_0_46# a_544_n15# a_0_94# VDD sky130_fd_pr__pfet_01v8 w=240 l=15
+  ad=7200 pd=540 as=6960 ps=665.6
XM1007 a_444_n15# a_344_n15# a_0_n15# GND sky130_fd_pr__nfet_01v8 w=42 l=15
+  ad=1218 pd=142 as=1218 ps=124.6
XM1008 a_544_n15# a_444_n15# a_0_n15# GND sky130_fd_pr__nfet_01v8 w=42 l=15
+  ad=1218 pd=142 as=1218 ps=124.6
XM1009 Clk_Out a_0_46# VDD VDD sky130_fd_pr__pfet_01v8 w=108 l=15
+  ad=3132 pd=274 as=3132 ps=278.64
XM1010 a_344_n15# a_244_n15# a_0_n15# GND sky130_fd_pr__nfet_01v8 w=42 l=15
+  ad=1218 pd=142 as=1218 ps=124.6
XM1011 a_544_n15# a_444_n15# a_0_94# VDD sky130_fd_pr__pfet_01v8 w=42 l=15
+  ad=1218 pd=142 as=1218 ps=116.48
XM1012 a_144_n15# a_44_n15# a_0_n15# GND sky130_fd_pr__nfet_01v8 w=42 l=15
+  ad=1218 pd=142 as=1218 ps=124.6
XM1013 a_244_n15# a_144_n15# a_0_n15# GND sky130_fd_pr__nfet_01v8 w=42 l=15
+  ad=1218 pd=142 as=1218 ps=124.6
XM1014 a_444_n15# a_344_n15# a_0_94# VDD sky130_fd_pr__pfet_01v8 w=42 l=15
+  ad=1218 pd=142 as=1218 ps=116.48
XM1015 a_44_n15# a_0_46# a_0_n15# GND sky130_fd_pr__nfet_01v8 w=42 l=15
+  ad=1218 pd=142 as=1218 ps=124.6
XM1016 a_344_n15# a_244_n15# a_0_94# VDD sky130_fd_pr__pfet_01v8 w=42 l=15
+  ad=1218 pd=142 as=1218 ps=116.48
XM1017 GND VCtrl a_n90_303# GND sky130_fd_pr__nfet_01v8 w=84 l=15
+  ad=2436 pd=227.415 as=2436 ps=226
XM1018 VDD a_n90_303# a_n90_303# VDD sky130_fd_pr__pfet_01v8 w=84 l=15
+  ad=2436 pd=216.72 as=2436 ps=226
XM1019 a_244_n15# a_144_n15# a_0_94# VDD sky130_fd_pr__pfet_01v8 w=42 l=15
+  ad=1218 pd=142 as=1218 ps=116.48
C0 a_0_n15# GND 2.20fF


v1 VDD 0 1.8
v2 VCtrl 0 0.8

.ic v(Clk_Out) = 0
.control 
tran 1ns 5us
plot v(Clk_Out)
.endc
