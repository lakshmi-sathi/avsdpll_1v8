magic
tech sky130A
timestamp 1606010604
<< nwell >>
rect 2951 1090 3441 1091
rect 2942 981 3441 1090
rect 3071 876 3118 981
rect 1033 856 1145 857
rect 2069 856 2116 857
rect 1033 847 1388 856
rect 862 799 1388 847
rect 1573 799 1660 856
rect 1845 800 2116 856
rect 2118 810 2162 869
rect 1845 799 2627 800
rect 862 698 2627 799
rect 862 670 2642 698
rect 847 669 2642 670
rect 847 659 891 669
rect 867 575 891 659
rect 1040 668 2627 669
rect 1040 642 2619 668
rect 867 571 904 575
rect 867 552 910 571
rect 867 526 961 552
rect 867 525 910 526
rect 867 506 891 525
rect 855 214 893 354
rect 809 78 945 214
<< locali >>
rect 2018 1294 2035 1311
rect 2052 1294 2069 1311
rect 2086 1294 2103 1311
rect 2030 1177 2068 1185
rect 2030 1174 2069 1177
rect 928 1157 965 1170
rect 928 1140 932 1157
rect 949 1140 965 1157
rect 2030 1157 2042 1174
rect 2059 1157 2069 1174
rect 2030 1154 2069 1157
rect 928 1131 965 1140
rect 1851 1137 2076 1154
rect 2021 1118 2076 1137
rect 2021 1094 2121 1118
rect 1944 1081 1979 1084
rect 1944 1064 1948 1081
rect 1965 1064 1979 1081
rect 1944 1055 1979 1064
rect 1944 1038 2114 1055
rect 54 852 129 880
rect 2097 875 2114 1038
rect 3015 911 3051 913
rect 3015 907 3019 911
rect 3007 887 3019 907
rect 3015 886 3019 887
rect 3048 886 3051 911
rect 3015 884 3051 886
rect 54 275 82 852
rect 1023 834 1056 875
rect 2058 858 2114 875
rect 1023 817 1161 834
rect 847 659 870 670
rect 874 552 910 561
rect 874 551 961 552
rect 874 534 877 551
rect 894 534 961 551
rect 874 526 961 534
rect 874 525 910 526
rect 740 490 777 498
rect 740 473 756 490
rect 773 473 777 490
rect 740 465 777 473
rect 2907 434 2995 448
rect 2907 417 2958 434
rect 2975 417 2995 434
rect 2907 394 2995 417
rect 863 370 885 375
rect 39 270 82 275
rect 39 248 45 270
rect 76 248 82 270
rect 39 244 82 248
rect 871 234 901 237
rect 871 217 878 234
rect 895 217 901 234
rect 871 205 901 217
rect 157 194 194 195
rect 157 184 195 194
rect 157 167 168 184
rect 185 167 195 184
rect 766 175 901 205
rect 157 157 195 167
rect 847 75 868 78
<< viali >>
rect 2035 1294 2052 1311
rect 2069 1294 2086 1311
rect 2103 1294 2120 1311
rect 932 1140 949 1157
rect 2042 1157 2059 1174
rect 1948 1064 1965 1081
rect 3019 886 3048 911
rect 877 534 894 551
rect 756 473 773 490
rect 2958 417 2975 434
rect 45 248 76 270
rect 878 217 895 234
rect 168 167 185 184
<< metal1 >>
rect 1842 1311 2163 1327
rect 1842 1294 2035 1311
rect 2052 1294 2069 1311
rect 2086 1294 2103 1311
rect 2120 1294 2163 1311
rect 1842 1278 2163 1294
rect 2991 1278 3217 1326
rect 2034 1179 2066 1182
rect 923 1163 958 1166
rect 923 1135 926 1163
rect 954 1135 958 1163
rect 2034 1153 2037 1179
rect 2063 1153 2066 1179
rect 2034 1150 2066 1153
rect 3138 1165 3217 1278
rect 3138 1164 3560 1165
rect 923 1132 958 1135
rect 3138 1124 3562 1164
rect 3138 1123 3513 1124
rect 1940 1086 1972 1089
rect 1940 1060 1943 1086
rect 1969 1060 1972 1086
rect 1940 1057 1972 1060
rect 0 975 31 989
rect 59 975 125 1006
rect 0 958 125 975
rect 3528 996 3562 1124
rect 3587 996 3618 1018
rect 3448 965 3502 966
rect 0 912 90 958
rect 3448 939 3473 965
rect 3499 939 3502 965
rect 3448 937 3502 939
rect 3528 934 3618 996
rect 3587 927 3618 934
rect 0 898 31 912
rect 3005 911 3053 919
rect 3005 886 3019 911
rect 3048 886 3053 911
rect 3005 877 3053 886
rect 3521 881 3553 882
rect 3443 879 3553 881
rect 2136 841 2180 869
rect 3443 853 3524 879
rect 3550 853 3553 879
rect 3443 851 3553 853
rect 3521 850 3553 851
rect 2136 815 2141 841
rect 2167 815 2180 841
rect 2136 810 2180 815
rect 0 734 31 741
rect 0 667 123 734
rect 1143 671 2925 703
rect 0 650 32 667
rect 101 639 123 667
rect 847 659 870 670
rect 2614 668 2627 671
rect 869 557 904 561
rect 869 528 872 557
rect 901 528 904 557
rect 869 525 904 528
rect 745 497 785 501
rect 0 466 31 483
rect 745 467 749 497
rect 780 467 785 497
rect 0 423 102 466
rect 745 463 785 467
rect 0 392 31 423
rect 65 390 102 423
rect 2951 439 2983 442
rect 2951 413 2954 439
rect 2980 413 2983 439
rect 2951 410 2983 413
rect 65 342 166 390
rect 863 370 885 375
rect 39 274 173 275
rect 39 270 199 274
rect 39 248 45 270
rect 76 248 199 270
rect 39 247 199 248
rect 39 244 82 247
rect 870 240 903 243
rect 870 212 873 240
rect 900 212 903 240
rect 870 209 903 212
rect 160 189 192 192
rect 160 163 163 189
rect 189 163 192 189
rect 160 160 192 163
rect 847 75 868 78
rect 2853 54 2904 55
rect 2775 46 2904 54
rect 2853 31 2904 46
rect 2832 0 2923 31
<< via1 >>
rect 926 1157 954 1163
rect 926 1140 932 1157
rect 932 1140 949 1157
rect 949 1140 954 1157
rect 926 1135 954 1140
rect 2037 1174 2063 1179
rect 2037 1157 2042 1174
rect 2042 1157 2059 1174
rect 2059 1157 2063 1174
rect 2037 1153 2063 1157
rect 1943 1081 1969 1086
rect 1943 1064 1948 1081
rect 1948 1064 1965 1081
rect 1965 1064 1969 1081
rect 1943 1060 1969 1064
rect 3473 939 3499 965
rect 3524 853 3550 879
rect 2141 815 2167 841
rect 872 551 901 557
rect 872 534 877 551
rect 877 534 894 551
rect 894 534 901 551
rect 872 528 901 534
rect 749 490 780 497
rect 749 473 756 490
rect 756 473 773 490
rect 773 473 780 490
rect 749 467 780 473
rect 2954 434 2980 439
rect 2954 417 2958 434
rect 2958 417 2975 434
rect 2975 417 2980 434
rect 2954 413 2980 417
rect 873 234 900 240
rect 873 217 878 234
rect 878 217 895 234
rect 895 217 900 234
rect 873 212 900 217
rect 163 184 189 189
rect 163 167 168 184
rect 168 167 185 184
rect 185 167 189 184
rect 163 163 189 167
<< metal2 >>
rect 1918 1343 1995 1371
rect 1942 1278 1970 1343
rect 1937 1273 1975 1278
rect 1937 1245 1942 1273
rect 1970 1245 1975 1273
rect 1937 1241 1975 1245
rect 2031 1180 2069 1185
rect 921 1163 960 1168
rect 921 1134 926 1163
rect 954 1134 960 1163
rect 2031 1152 2036 1180
rect 2064 1152 2069 1180
rect 2031 1147 2069 1152
rect 921 1129 960 1134
rect 1937 1087 1975 1092
rect 1937 1059 1942 1087
rect 1970 1059 1975 1087
rect 1937 1054 1975 1059
rect 289 1020 1974 1021
rect 289 992 2172 1020
rect 0 828 28 854
rect 289 828 320 992
rect 1804 991 2172 992
rect 2138 846 2172 991
rect 3470 965 3502 966
rect 3470 939 3473 965
rect 3499 939 3502 965
rect 3182 870 3208 894
rect 0 799 320 828
rect 2136 841 2172 846
rect 2136 815 2141 841
rect 2167 815 2172 841
rect 2136 809 2172 815
rect 0 777 28 799
rect 3259 765 3261 789
rect 3259 745 3287 765
rect 2872 715 3289 745
rect 2872 703 2925 715
rect 302 671 2925 703
rect 3470 686 3502 939
rect 3590 882 3618 904
rect 3521 879 3618 882
rect 3521 853 3524 879
rect 3550 853 3618 879
rect 3521 850 3618 853
rect 3590 827 3618 850
rect 0 584 28 606
rect 302 584 335 671
rect 0 552 335 584
rect 869 557 904 671
rect 0 529 28 552
rect 869 528 872 557
rect 901 528 904 557
rect 869 525 904 528
rect 3032 654 3502 686
rect 745 497 785 501
rect 745 467 749 497
rect 780 467 785 497
rect 745 370 785 467
rect 3032 442 3067 654
rect 2951 439 3067 442
rect 2951 413 2954 439
rect 2980 413 3067 439
rect 2951 410 3067 413
rect 694 330 785 370
rect 157 190 195 195
rect 157 162 162 190
rect 190 162 195 190
rect 157 157 195 162
rect 694 144 734 330
rect 870 240 903 318
rect 870 212 873 240
rect 900 212 903 240
rect 870 209 903 212
rect 2919 186 2992 192
rect 868 144 909 155
rect 694 104 909 144
rect 2919 120 2925 186
rect 2985 157 2992 186
rect 2985 120 3034 157
rect 2919 114 3034 120
rect 2981 28 3034 114
rect 2969 0 3046 28
<< via2 >>
rect 1942 1245 1970 1273
rect 926 1135 954 1162
rect 926 1134 954 1135
rect 2036 1179 2064 1180
rect 2036 1153 2037 1179
rect 2037 1153 2063 1179
rect 2063 1153 2064 1179
rect 2036 1152 2064 1153
rect 1942 1086 1970 1087
rect 1942 1060 1943 1086
rect 1943 1060 1969 1086
rect 1969 1060 1970 1086
rect 1942 1059 1970 1060
rect 162 189 190 190
rect 162 163 163 189
rect 163 163 189 189
rect 189 163 190 189
rect 162 162 190 163
rect 2925 120 2985 186
<< metal3 >>
rect 725 1273 1979 1282
rect 725 1245 1942 1273
rect 1970 1245 1979 1273
rect 725 1244 1979 1245
rect 725 1097 763 1244
rect 1934 1236 1979 1244
rect 2031 1180 2093 1185
rect 891 1162 960 1168
rect 891 1134 926 1162
rect 954 1134 960 1162
rect 2031 1152 2036 1180
rect 2064 1157 2093 1180
rect 2064 1152 2094 1157
rect 2031 1147 2094 1152
rect 891 1129 960 1134
rect 725 998 764 1097
rect 891 1061 926 1129
rect 1937 1087 1975 1092
rect 1937 1061 1942 1087
rect 891 1059 1942 1061
rect 1970 1085 1975 1087
rect 1970 1059 1979 1085
rect 891 1026 1979 1059
rect 501 987 764 998
rect 501 960 763 987
rect 501 435 539 960
rect 2055 555 2094 1147
rect 2055 554 2293 555
rect 2055 514 2330 554
rect 337 397 539 435
rect 2268 437 2330 514
rect 337 195 375 397
rect 2268 230 2331 437
rect 157 190 375 195
rect 157 162 162 190
rect 190 162 375 190
rect 157 157 375 162
rect 2269 161 2331 230
rect 2919 186 2992 192
rect 2919 161 2925 186
rect 2269 120 2925 161
rect 2985 120 2992 186
rect 2269 113 2992 120
use FD  FD_2
timestamp 1605926473
transform -1 0 1867 0 1 1006
box 0 0 935 320
use FD  FD_0
timestamp 1605926473
transform -1 0 1034 0 -1 1006
box 0 0 935 320
use PFD  PFD_0
timestamp 1605977318
transform 1 0 101 0 1 46
box 0 0 767 640
use FD  FD_1
timestamp 1605926473
transform -1 0 2075 0 -1 1006
box 0 0 935 320
use CP  CP_0
timestamp 1605998167
transform 1 0 867 0 1 46
box 0 0 2067 640
use VCO  VCO_0
timestamp 1605977318
transform -1 0 3016 0 -1 1326
box 0 0 902 640
use MUX  MUX_0
timestamp 1605906497
transform -1 0 3453 0 1 743
box 0 -12 408 285
<< labels >>
rlabel metal1 2832 0 2923 0 1 VDD#2
port 7 n power bidirectional
rlabel metal2 2969 0 3046 0 1 CLK
port 4 n signal output
rlabel metal2 1918 1371 1995 1371 5 REF
port 10 s signal input
rlabel metal1 3618 927 3618 1018 7 VDD#3
port 9 w power bidirectional
rlabel metal2 3618 827 3618 904 7 VCO_IN
port 8 w signal input
rlabel metal1 0 392 0 483 3 GND#2
port 6 e ground bidirectional
rlabel metal2 0 777 0 854 3 ENb_VCO
port 5 e signal input
rlabel metal2 0 529 0 606 3 ENb_CP
port 3 e signal input
rlabel metal1 0 650 0 741 3 VDD
port 2 e power bidirectional
rlabel metal1 0 898 0 989 3 GND
port 1 e ground bidirectional
<< properties >>
string LEFclass CORE
string LEFsite unithddb1
<< end >>
