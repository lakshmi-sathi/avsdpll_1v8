magic
tech sky130A
timestamp 1605147420
<< nwell >>
rect -103 429 793 514
rect 265 185 793 429
rect -61 76 793 185
<< nmos >>
rect -61 303 -46 387
rect 10 249 118 264
rect 29 -15 44 27
rect 129 -15 144 27
rect 229 -15 244 27
rect 329 -15 344 27
rect 429 -15 444 27
rect 529 -15 544 27
rect 629 -93 644 27
rect 731 -26 746 28
<< pmos >>
rect 461 302 476 386
rect 284 244 392 259
rect 29 94 44 136
rect 129 94 144 136
rect 229 94 244 136
rect 329 94 344 136
rect 429 94 444 136
rect 529 94 544 136
rect 629 94 644 334
rect 731 94 746 202
<< ndiff >>
rect -90 365 -61 387
rect -90 347 -84 365
rect -67 347 -61 365
rect -90 329 -61 347
rect -90 311 -84 329
rect -67 311 -61 329
rect -90 303 -61 311
rect -46 364 -17 387
rect -46 347 -40 364
rect -23 347 -17 364
rect -46 329 -17 347
rect -46 311 -40 329
rect -23 311 -17 329
rect -46 303 -17 311
rect 10 287 118 293
rect 10 270 18 287
rect 35 270 52 287
rect 69 270 86 287
rect 103 270 118 287
rect 10 264 118 270
rect 10 243 118 249
rect 10 226 14 243
rect 31 226 48 243
rect 65 226 82 243
rect 99 226 118 243
rect 10 220 118 226
rect 0 14 29 27
rect 0 -3 6 14
rect 23 -3 29 14
rect 0 -15 29 -3
rect 44 14 73 27
rect 44 -3 50 14
rect 67 -3 73 14
rect 44 -15 73 -3
rect 100 14 129 27
rect 100 -3 106 14
rect 123 -3 129 14
rect 100 -15 129 -3
rect 144 14 173 27
rect 144 -3 150 14
rect 167 -3 173 14
rect 144 -15 173 -3
rect 200 14 229 27
rect 200 -3 206 14
rect 223 -3 229 14
rect 200 -15 229 -3
rect 244 14 273 27
rect 244 -3 250 14
rect 267 -3 273 14
rect 244 -15 273 -3
rect 300 14 329 27
rect 300 -3 306 14
rect 323 -3 329 14
rect 300 -15 329 -3
rect 344 14 373 27
rect 344 -3 350 14
rect 367 -3 373 14
rect 344 -15 373 -3
rect 400 14 429 27
rect 400 -3 406 14
rect 423 -3 429 14
rect 400 -15 429 -3
rect 444 14 473 27
rect 444 -3 450 14
rect 467 -3 473 14
rect 444 -15 473 -3
rect 500 14 529 27
rect 500 -3 506 14
rect 523 -3 529 14
rect 500 -15 529 -3
rect 544 14 573 27
rect 544 -3 550 14
rect 567 -3 573 14
rect 544 -15 573 -3
rect 600 14 629 27
rect 600 -3 606 14
rect 623 -3 629 14
rect 600 -20 629 -3
rect 600 -37 606 -20
rect 623 -37 629 -20
rect 600 -54 629 -37
rect 600 -71 606 -54
rect 623 -71 629 -54
rect 600 -93 629 -71
rect 644 14 673 27
rect 644 -3 650 14
rect 667 -3 673 14
rect 644 -20 673 -3
rect 644 -37 650 -20
rect 667 -37 673 -20
rect 702 8 731 28
rect 702 -9 708 8
rect 725 -9 731 8
rect 702 -26 731 -9
rect 746 8 775 28
rect 746 -9 752 8
rect 769 -9 775 8
rect 746 -26 775 -9
rect 644 -54 673 -37
rect 644 -71 650 -54
rect 667 -71 673 -54
rect 644 -93 673 -71
<< pdiff >>
rect 432 378 461 386
rect 432 361 438 378
rect 455 361 461 378
rect 432 344 461 361
rect 432 327 438 344
rect 455 327 461 344
rect 432 302 461 327
rect 476 382 505 386
rect 476 365 482 382
rect 499 365 505 382
rect 476 348 505 365
rect 476 331 482 348
rect 499 331 505 348
rect 476 302 505 331
rect 284 282 392 288
rect 284 265 292 282
rect 309 265 326 282
rect 343 265 360 282
rect 377 265 392 282
rect 284 259 392 265
rect 600 292 629 334
rect 600 275 606 292
rect 623 275 629 292
rect 600 250 629 275
rect 284 238 392 244
rect 284 221 292 238
rect 309 221 326 238
rect 343 221 360 238
rect 377 221 392 238
rect 284 215 392 221
rect 600 233 606 250
rect 623 233 629 250
rect 600 208 629 233
rect 600 191 606 208
rect 623 191 629 208
rect 600 166 629 191
rect 600 149 606 166
rect 623 149 629 166
rect 0 124 29 136
rect 0 107 6 124
rect 23 107 29 124
rect 0 94 29 107
rect 44 124 73 136
rect 44 107 50 124
rect 67 107 73 124
rect 44 94 73 107
rect 100 124 129 136
rect 100 107 106 124
rect 123 107 129 124
rect 100 94 129 107
rect 144 124 173 136
rect 144 107 150 124
rect 167 107 173 124
rect 144 94 173 107
rect 200 124 229 136
rect 200 107 206 124
rect 223 107 229 124
rect 200 94 229 107
rect 244 124 273 136
rect 244 107 250 124
rect 267 107 273 124
rect 244 94 273 107
rect 300 124 329 136
rect 300 107 306 124
rect 323 107 329 124
rect 300 94 329 107
rect 344 124 373 136
rect 344 107 350 124
rect 367 107 373 124
rect 344 94 373 107
rect 400 124 429 136
rect 400 107 406 124
rect 423 107 429 124
rect 400 94 429 107
rect 444 124 473 136
rect 444 107 450 124
rect 467 107 473 124
rect 444 94 473 107
rect 500 124 529 136
rect 500 107 506 124
rect 523 107 529 124
rect 500 94 529 107
rect 544 124 573 136
rect 544 107 550 124
rect 567 107 573 124
rect 544 94 573 107
rect 600 124 629 149
rect 600 107 606 124
rect 623 107 629 124
rect 600 94 629 107
rect 644 292 674 334
rect 644 275 650 292
rect 667 275 674 292
rect 644 250 674 275
rect 644 233 650 250
rect 667 233 674 250
rect 644 208 674 233
rect 644 191 650 208
rect 667 191 674 208
rect 644 166 674 191
rect 644 149 650 166
rect 667 149 674 166
rect 644 124 674 149
rect 644 107 650 124
rect 667 107 674 124
rect 644 94 674 107
rect 702 196 731 202
rect 702 178 708 196
rect 725 178 731 196
rect 702 160 731 178
rect 702 142 708 160
rect 725 142 731 160
rect 702 124 731 142
rect 702 107 708 124
rect 725 107 731 124
rect 702 94 731 107
rect 746 189 775 202
rect 746 172 752 189
rect 769 172 775 189
rect 746 154 775 172
rect 746 136 752 154
rect 769 136 775 154
rect 746 118 775 136
rect 746 100 752 118
rect 769 100 775 118
rect 746 94 775 100
<< ndiffc >>
rect -84 347 -67 365
rect -84 311 -67 329
rect -40 347 -23 364
rect -40 311 -23 329
rect 18 270 35 287
rect 52 270 69 287
rect 86 270 103 287
rect 14 226 31 243
rect 48 226 65 243
rect 82 226 99 243
rect 6 -3 23 14
rect 50 -3 67 14
rect 106 -3 123 14
rect 150 -3 167 14
rect 206 -3 223 14
rect 250 -3 267 14
rect 306 -3 323 14
rect 350 -3 367 14
rect 406 -3 423 14
rect 450 -3 467 14
rect 506 -3 523 14
rect 550 -3 567 14
rect 606 -3 623 14
rect 606 -37 623 -20
rect 606 -71 623 -54
rect 650 -3 667 14
rect 650 -37 667 -20
rect 708 -9 725 8
rect 752 -9 769 8
rect 650 -71 667 -54
<< pdiffc >>
rect 438 361 455 378
rect 438 327 455 344
rect 482 365 499 382
rect 482 331 499 348
rect 292 265 309 282
rect 326 265 343 282
rect 360 265 377 282
rect 606 275 623 292
rect 292 221 309 238
rect 326 221 343 238
rect 360 221 377 238
rect 606 233 623 250
rect 606 191 623 208
rect 606 149 623 166
rect 6 107 23 124
rect 50 107 67 124
rect 106 107 123 124
rect 150 107 167 124
rect 206 107 223 124
rect 250 107 267 124
rect 306 107 323 124
rect 350 107 367 124
rect 406 107 423 124
rect 450 107 467 124
rect 506 107 523 124
rect 550 107 567 124
rect 606 107 623 124
rect 650 275 667 292
rect 650 233 667 250
rect 650 191 667 208
rect 650 149 667 166
rect 650 107 667 124
rect 708 178 725 196
rect 708 142 725 160
rect 708 107 725 124
rect 752 172 769 189
rect 752 136 769 154
rect 752 100 769 118
<< psubdiff >>
rect 37 332 49 364
rect 81 332 93 364
rect 37 320 93 332
rect -90 -146 -78 -122
rect -54 -146 -42 -122
rect 6 -146 18 -122
rect 42 -146 54 -122
rect 102 -146 114 -122
rect 138 -146 150 -122
rect 198 -146 210 -122
rect 234 -146 246 -122
rect 294 -146 306 -122
rect 330 -146 342 -122
rect 390 -146 402 -122
rect 426 -146 438 -122
rect 486 -146 498 -122
rect 522 -146 534 -122
rect 582 -146 594 -122
rect 618 -146 630 -122
rect 678 -146 690 -122
rect 714 -146 726 -122
<< nsubdiff >>
rect -85 461 -73 485
rect -49 461 -37 485
rect 11 461 23 485
rect 47 461 59 485
rect 107 461 119 485
rect 143 461 155 485
rect 203 461 215 485
rect 239 461 251 485
rect 299 461 311 485
rect 335 461 347 485
rect 395 461 407 485
rect 431 461 443 485
rect 491 461 503 485
rect 527 461 539 485
rect 587 461 599 485
rect 623 461 635 485
rect 683 461 695 485
rect 719 461 731 485
<< psubdiffcont >>
rect 49 332 81 364
rect -78 -146 -54 -122
rect 18 -146 42 -122
rect 114 -146 138 -122
rect 210 -146 234 -122
rect 306 -146 330 -122
rect 402 -146 426 -122
rect 498 -146 522 -122
rect 594 -146 618 -122
rect 690 -146 714 -122
<< nsubdiffcont >>
rect -73 461 -49 485
rect 23 461 47 485
rect 119 461 143 485
rect 215 461 239 485
rect 311 461 335 485
rect 407 461 431 485
rect 503 461 527 485
rect 599 461 623 485
rect 695 461 719 485
<< poly >>
rect -61 387 -46 400
rect 352 396 476 416
rect 352 386 375 396
rect 461 386 476 396
rect 342 375 375 386
rect 342 358 350 375
rect 367 358 375 375
rect 342 353 375 358
rect -61 289 -46 303
rect 629 334 644 347
rect -61 288 -27 289
rect -62 278 -27 288
rect -62 261 -54 278
rect -37 264 -27 278
rect -37 261 10 264
rect -62 249 10 261
rect 118 249 131 264
rect 461 259 476 302
rect 271 244 284 259
rect 392 244 476 259
rect 29 136 44 149
rect 129 136 144 149
rect 229 136 244 149
rect 329 136 344 149
rect 429 136 444 149
rect 529 136 544 149
rect 731 202 746 215
rect 29 86 44 94
rect 129 86 144 94
rect 229 86 244 94
rect 329 86 344 94
rect 429 86 444 94
rect 529 86 544 94
rect 629 86 644 94
rect 22 76 44 86
rect 122 76 144 86
rect 222 76 244 86
rect 322 76 344 86
rect 422 76 444 86
rect 522 76 544 86
rect 622 76 644 86
rect 0 69 44 76
rect 0 52 8 69
rect 25 52 44 69
rect 0 46 44 52
rect 100 69 144 76
rect 100 52 108 69
rect 125 52 144 69
rect 100 46 144 52
rect 200 69 244 76
rect 200 52 208 69
rect 225 52 244 69
rect 200 46 244 52
rect 300 69 344 76
rect 300 52 308 69
rect 325 52 344 69
rect 300 46 344 52
rect 400 69 444 76
rect 400 52 408 69
rect 425 52 444 69
rect 400 46 444 52
rect 500 69 544 76
rect 500 52 508 69
rect 525 52 544 69
rect 500 46 544 52
rect 600 69 644 76
rect 731 75 746 94
rect 600 52 608 69
rect 625 52 644 69
rect 600 46 644 52
rect 701 69 746 75
rect 701 52 709 69
rect 726 52 746 69
rect 701 46 746 52
rect 22 35 44 46
rect 122 35 144 46
rect 222 35 244 46
rect 322 35 344 46
rect 422 35 444 46
rect 522 35 544 46
rect 622 35 644 46
rect 29 27 44 35
rect 129 27 144 35
rect 229 27 244 35
rect 329 27 344 35
rect 429 27 444 35
rect 529 27 544 35
rect 629 27 644 35
rect 731 28 746 46
rect 29 -28 44 -15
rect 129 -28 144 -15
rect 229 -28 244 -15
rect 329 -28 344 -15
rect 429 -28 444 -15
rect 529 -28 544 -15
rect 731 -39 746 -26
rect 629 -106 644 -93
<< polycont >>
rect 350 358 367 375
rect -54 261 -37 278
rect 8 52 25 69
rect 108 52 125 69
rect 208 52 225 69
rect 308 52 325 69
rect 408 52 425 69
rect 508 52 525 69
rect 608 52 625 69
rect 709 52 726 69
<< locali >>
rect -103 485 793 514
rect -103 461 -73 485
rect -49 461 23 485
rect 47 461 119 485
rect 143 461 215 485
rect 239 461 311 485
rect 335 461 407 485
rect 431 461 503 485
rect 527 461 599 485
rect 623 461 695 485
rect 719 461 793 485
rect -103 438 793 461
rect 478 437 510 438
rect -84 406 89 421
rect 482 414 510 437
rect -84 404 193 406
rect -84 365 -67 404
rect -84 329 -67 347
rect -84 303 -67 311
rect -40 364 -23 387
rect 30 386 193 404
rect 30 385 321 386
rect 145 377 321 385
rect 438 378 455 386
rect 145 375 375 377
rect 145 365 350 375
rect -23 347 49 364
rect -40 332 49 347
rect 81 332 100 364
rect 261 358 350 365
rect 367 366 375 375
rect 367 361 438 366
rect 367 358 455 361
rect 261 345 455 358
rect -40 329 100 332
rect -23 319 100 329
rect 363 344 455 345
rect 363 327 438 344
rect 363 325 455 327
rect -40 303 -23 311
rect 30 287 100 319
rect 438 302 455 325
rect 482 382 502 414
rect 499 365 502 382
rect 482 348 502 365
rect 499 331 502 348
rect 482 295 502 331
rect 708 354 749 438
rect -102 278 -29 280
rect -102 261 -54 278
rect -37 261 -29 278
rect 10 270 18 287
rect 35 270 52 287
rect 69 270 86 287
rect 103 270 118 287
rect 476 282 502 295
rect 284 265 292 282
rect 309 265 326 282
rect 343 265 360 282
rect 377 265 502 282
rect 606 292 623 317
rect -102 260 -29 261
rect 606 250 623 275
rect -88 226 14 243
rect 31 226 48 243
rect 65 226 82 243
rect 99 226 119 243
rect -88 218 119 226
rect 284 221 292 238
rect 309 221 326 238
rect 343 221 360 238
rect 377 221 392 238
rect 534 233 606 250
rect -88 -32 -51 218
rect 306 185 365 221
rect 534 215 623 233
rect 474 208 623 215
rect 474 191 606 208
rect 474 185 623 191
rect 6 166 623 185
rect 6 153 606 166
rect 6 124 23 153
rect 6 94 23 107
rect 50 124 67 136
rect 50 69 67 107
rect 106 124 123 153
rect 106 94 123 107
rect 150 124 167 136
rect 150 69 167 107
rect 206 124 223 153
rect 206 94 223 107
rect 250 124 267 136
rect 250 69 267 107
rect 306 124 323 153
rect 306 94 323 107
rect 350 124 367 136
rect 350 69 367 107
rect 406 124 423 153
rect 406 94 423 107
rect 450 124 467 136
rect 450 69 467 107
rect 506 124 523 153
rect 506 94 523 107
rect 550 124 567 136
rect 550 69 567 107
rect 606 124 623 149
rect 606 94 623 107
rect 650 292 667 317
rect 650 250 667 275
rect 650 208 667 233
rect 650 166 667 191
rect 650 124 667 149
rect 650 75 667 107
rect 708 281 738 354
rect 708 196 725 281
rect 708 160 725 178
rect 708 124 725 142
rect 708 94 725 107
rect 752 189 769 202
rect 752 154 769 172
rect 752 118 769 136
rect 650 69 734 75
rect -10 52 8 69
rect 25 52 33 69
rect 50 52 108 69
rect 125 52 133 69
rect 150 52 208 69
rect 225 52 233 69
rect 250 52 308 69
rect 325 52 333 69
rect 350 52 408 69
rect 425 52 433 69
rect 450 52 508 69
rect 525 52 533 69
rect 550 52 608 69
rect 625 52 633 69
rect 650 52 683 69
rect 700 52 709 69
rect 726 52 734 69
rect 6 14 23 27
rect 6 -32 23 -3
rect 50 14 67 52
rect 50 -15 67 -3
rect 106 14 123 27
rect 106 -32 123 -3
rect 150 14 167 52
rect 150 -15 167 -3
rect 206 14 223 27
rect 206 -32 223 -3
rect 250 14 267 52
rect 250 -15 267 -3
rect 306 14 323 27
rect 306 -32 323 -3
rect 350 14 367 52
rect 350 -15 367 -3
rect 406 14 423 27
rect 406 -32 423 -3
rect 450 14 467 52
rect 450 -15 467 -3
rect 506 14 523 27
rect 506 -32 523 -3
rect 550 14 567 52
rect 650 46 734 52
rect 752 72 769 100
rect 752 49 793 72
rect 550 -15 567 -3
rect 606 14 623 27
rect 606 -20 623 -3
rect 591 -32 606 -26
rect -88 -37 606 -32
rect -88 -54 623 -37
rect -88 -64 606 -54
rect 591 -69 606 -64
rect 606 -82 623 -71
rect 650 14 667 46
rect 650 -20 667 -3
rect 650 -54 667 -37
rect 708 8 725 28
rect 708 -43 725 -9
rect 752 8 769 49
rect 752 -26 769 -9
rect 650 -82 667 -71
rect 703 -74 726 -43
rect 699 -110 726 -74
rect -104 -122 795 -110
rect -104 -146 -78 -122
rect -54 -146 18 -122
rect 42 -146 114 -122
rect 138 -146 210 -122
rect 234 -146 306 -122
rect 330 -146 402 -122
rect 426 -146 498 -122
rect 522 -146 594 -122
rect 618 -146 690 -122
rect 714 -146 795 -122
rect -104 -158 795 -146
<< viali >>
rect -27 52 -10 69
rect 683 52 700 69
<< metal1 >>
rect -33 69 704 75
rect -33 52 -27 69
rect -10 52 683 69
rect 700 52 704 69
rect -33 47 704 52
rect -33 46 703 47
<< labels >>
rlabel locali -102 260 -102 280 3 VCtrl
port 2 e
rlabel locali -103 438 -103 514 3 VDD
port 3 e
rlabel locali -104 -158 -104 -110 3 GND
port 1 e
rlabel locali 793 49 793 72 7 Clk_Out
port 4 w
<< end >>
